-- megafunction wizard: %ALTFP_DIV%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altfp_div 

-- ============================================================
-- File Name: k_ukf_div.vhd
-- Megafunction Name(s):
-- 			altfp_div
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.1 Build 259 01/25/2012 SP 2 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altfp_div CBX_AUTO_BLACKBOX="ALL" DENORMAL_SUPPORT="NO" DEVICE_FAMILY="Cyclone II" OPTIMIZE="SPEED" PIPELINE=14 REDUCED_FUNCTIONALITY="NO" WIDTH_EXP=8 WIDTH_MAN=23 clock dataa datab result
--VERSION_BEGIN 11.1SP2 cbx_altbarrel_shift 2012:01:25:21:13:53:SJ cbx_altfp_div 2012:01:25:21:13:53:SJ cbx_altsyncram 2012:01:25:21:13:53:SJ cbx_cycloneii 2012:01:25:21:13:53:SJ cbx_lpm_abs 2012:01:25:21:13:53:SJ cbx_lpm_add_sub 2012:01:25:21:13:53:SJ cbx_lpm_compare 2012:01:25:21:13:53:SJ cbx_lpm_decode 2012:01:25:21:13:53:SJ cbx_lpm_divide 2012:01:25:21:13:53:SJ cbx_lpm_mult 2012:01:25:21:13:53:SJ cbx_lpm_mux 2012:01:25:21:13:53:SJ cbx_mgl 2012:01:25:21:15:41:SJ cbx_padd 2012:01:25:21:13:53:SJ cbx_stratix 2012:01:25:21:13:53:SJ cbx_stratixii 2012:01:25:21:13:53:SJ cbx_stratixiii 2012:01:25:21:13:53:SJ cbx_stratixv 2012:01:25:21:13:53:SJ cbx_util_mgl 2012:01:25:21:13:53:SJ  VERSION_END


--altfp_div_pst CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" FILE_NAME="k_ukf_div.vhd:a" PIPELINE=14 WIDTH_EXP=8 WIDTH_MAN=23 aclr clk_en clock dataa datab result
--VERSION_BEGIN 11.1SP2 cbx_altbarrel_shift 2012:01:25:21:13:53:SJ cbx_altfp_div 2012:01:25:21:13:53:SJ cbx_altsyncram 2012:01:25:21:13:53:SJ cbx_cycloneii 2012:01:25:21:13:53:SJ cbx_lpm_abs 2012:01:25:21:13:53:SJ cbx_lpm_add_sub 2012:01:25:21:13:53:SJ cbx_lpm_compare 2012:01:25:21:13:53:SJ cbx_lpm_decode 2012:01:25:21:13:53:SJ cbx_lpm_divide 2012:01:25:21:13:53:SJ cbx_lpm_mult 2012:01:25:21:13:53:SJ cbx_lpm_mux 2012:01:25:21:13:53:SJ cbx_mgl 2012:01:25:21:15:41:SJ cbx_padd 2012:01:25:21:13:53:SJ cbx_stratix 2012:01:25:21:13:53:SJ cbx_stratixii 2012:01:25:21:13:53:SJ cbx_stratixiii 2012:01:25:21:13:53:SJ cbx_stratixv 2012:01:25:21:13:53:SJ cbx_util_mgl 2012:01:25:21:13:53:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = altsyncram 1 lpm_add_sub 4 lpm_compare 1 lpm_mult 5 mux21 74 reg 847 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  k_ukf_div_altfp_div_pst_o3f IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 datab	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END k_ukf_div_altfp_div_pst_o3f;

 ARCHITECTURE RTL OF k_ukf_div_altfp_div_pst_o3f IS

	 SIGNAL  wire_altsyncram3_q_a	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL	 a_is_infinity_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_is_infinity_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_a_is_infinity_dffe_1_w_lg_q318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 a_is_infinity_dffe_10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_is_infinity_dffe_11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_is_infinity_dffe_12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_is_infinity_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_is_infinity_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_is_infinity_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_is_infinity_dffe_5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_is_infinity_dffe_6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_is_infinity_dffe_7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_is_infinity_dffe_8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_is_infinity_dffe_9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_a_zero_b_not_dffe_1_w_lg_q326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 a_zero_b_not_dffe_10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b1_dffe_0	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b1_dffe_1	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_b_is_infinity_dffe_1_w_lg_q325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 b_is_infinity_dffe_10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 both_exp_zeros_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_divbyzero_pipe_dffe_1_w_lg_q317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 divbyzero_pipe_dffe_10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 e1_dffe_0	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 e1_dffe_1	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 e1_dffe_perf_0	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 e1_dffe_perf_1	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 e1_dffe_perf_2	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 e1_dffe_perf_3	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_0	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_1	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_10	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_11	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_2	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_3	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_4	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_5	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_6	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_7	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_8	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_9	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 frac_a_smaller_dffe1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_a_dffe1_dffe1	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_b_dffe1_dffe1	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_result_dffe	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_nan_pipe_dffe_1_w_lg_q308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 nan_pipe_dffe_10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 over_under_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 over_under_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 over_under_dffe_10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 over_under_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 over_under_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 over_under_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 over_under_dffe_5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 over_under_dffe_6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 over_under_dffe_7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 over_under_dffe_8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 over_under_dffe_9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_partial_perf_dffe_0	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_q_partial_perf_dffe_0_w_q_range373w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL	 q_partial_perf_dffe_1	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_q_partial_perf_dffe_1_w_lg_w_q_range407w408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_q_partial_perf_dffe_1_w_lg_w_q_range410w411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_q_partial_perf_dffe_1_w_lg_w_q_range413w414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_q_partial_perf_dffe_1_w_lg_w_q_range416w417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_q_partial_perf_dffe_1_w_q_range407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_q_partial_perf_dffe_1_w_q_range410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_q_partial_perf_dffe_1_w_q_range413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_q_partial_perf_dffe_1_w_q_range416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 quotient_j_dffe	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 quotient_k_dffe_0	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 quotient_k_dffe_perf_0	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 quotient_k_dffe_perf_1	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 quotient_k_dffe_perf_2	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 quotient_k_dffe_perf_3	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 remainder_j_dffe_0	:	STD_LOGIC_VECTOR(49 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 remainder_j_dffe_1	:	STD_LOGIC_VECTOR(49 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 remainder_j_dffe_perf_0	:	STD_LOGIC_VECTOR(49 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 remainder_j_dffe_perf_1	:	STD_LOGIC_VECTOR(49 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 remainder_j_dffe_perf_2	:	STD_LOGIC_VECTOR(49 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_bias_addition_overflow	:	STD_LOGIC;
	 SIGNAL  wire_bias_addition_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exp_sub_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_quotient_process_dataa	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_quotient_process_datab	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_quotient_process_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_quotient_process_w_result_range425w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_remainder_sub_0_dataa	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_remainder_sub_0_result	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_cmpr2_alb	:	STD_LOGIC;
	 SIGNAL  wire_a1_prod_datab	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_a1_prod_result	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  wire_b1_prod_w_lg_w_result_range359w360w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_b1_prod_datab	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_b1_prod_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_b1_prod_w_result_range359w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_q_partial_0_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_q_partial_1_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_remainder_mult_0_result	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL	wire_exp_result_muxa_dataout	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	wire_man_a_adjusteda_dataout	:	STD_LOGIC_VECTOR(24 DOWNTO 0);
	 SIGNAL	wire_man_result_muxa_dataout	:	STD_LOGIC_VECTOR(22 DOWNTO 0);
	 SIGNAL	wire_select_bias_2a_dataout	:	STD_LOGIC_VECTOR(8 DOWNTO 0);
	 SIGNAL	wire_select_biasa_dataout	:	STD_LOGIC_VECTOR(8 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_lg_w_lg_bias_addition_overf_w304w305w306w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w304w305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w304w312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w302w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range262w286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range265w288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range268w290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range271w292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range274w294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range277w296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range280w298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range11w18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range21w28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range31w38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range41w48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range51w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range61w68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range71w78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range14w20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range24w30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range34w40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range44w50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range54w60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range64w70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range74w80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_exp_a_all_one_w_range77w222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_exp_add_output_all_one_range297w321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_exp_b_all_one_w_range79w224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_exp_b_not_zero_w_range75w256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_a_is_infinity_w233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_a_is_nan_w234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_bias_addition_overf_w304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_exp_sign_w303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_exp_a_not_zero_w_range72w227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_man_a_not_zero_w_range214w221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_man_b_not_zero_w_range217w223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_lg_w_lg_bias_addition_overf_w299w300w301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w299w300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_bias_addition_overf_w323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_bias_addition_overf_w299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range262w264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range265w267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range268w270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range271w273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range274w276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range277w279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range280w282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range141w143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range147w149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range153w155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range159w161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range165w167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range171w173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range177w179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range183w185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range189w191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range195w197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range87w89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range201w203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range207w209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range213w215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range11w13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range21w23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range31w33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range41w43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range51w53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range61w63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range93w95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range71w73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range99w101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range105w107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range111w113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range117w119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range123w125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range129w131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range135w137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range144w146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range150w152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range156w158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range162w164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range168w170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range174w176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range180w182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range186w188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range192w194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range198w200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range90w92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range204w206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range210w212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range216w218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range14w16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range24w26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range34w36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range44w46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range54w56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range64w66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range96w98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range74w76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range102w104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range108w110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range114w116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range120w122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range126w128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range132w134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range138w140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  a_is_infinity_w :	STD_LOGIC;
	 SIGNAL  a_is_nan_w :	STD_LOGIC;
	 SIGNAL  a_zero_b_not :	STD_LOGIC;
	 SIGNAL  b1_dffe_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  b_is_infinity_w :	STD_LOGIC;
	 SIGNAL  b_is_nan_w :	STD_LOGIC;
	 SIGNAL  bias_addition_overf_w :	STD_LOGIC;
	 SIGNAL  bias_addition_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  both_exp_zeros :	STD_LOGIC;
	 SIGNAL  e0_dffe1_wo :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  e0_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  e1_w :	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  exp_a_all_one_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_a_not_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_add_output_all_one :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_add_output_not_zero :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_b_all_one_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_b_not_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_result_mux_out :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_result_mux_sel_w :	STD_LOGIC;
	 SIGNAL  exp_result_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_sign_w :	STD_LOGIC;
	 SIGNAL  exp_sub_a_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_sub_b_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_sub_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  frac_a_smaller_dffe1_wi :	STD_LOGIC;
	 SIGNAL  frac_a_smaller_dffe1_wo :	STD_LOGIC;
	 SIGNAL  frac_a_smaller_w :	STD_LOGIC;
	 SIGNAL  guard_bit :	STD_LOGIC;
	 SIGNAL  man_a_adjusted_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  man_a_dffe1_wi :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_a_dffe1_wo :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_a_not_zero_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_b_adjusted_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_b_dffe1_wi :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_b_dffe1_wo :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_b_not_zero_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_result_dffe_wi :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_result_dffe_wo :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_result_mux_select :	STD_LOGIC;
	 SIGNAL  man_result_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_zeros_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  overflow_ones_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  overflow_underflow :	STD_LOGIC;
	 SIGNAL  overflow_w :	STD_LOGIC;
	 SIGNAL  quotient_accumulate_w :	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  quotient_process_cin_w :	STD_LOGIC;
	 SIGNAL  remainder_j_w :	STD_LOGIC_VECTOR (99 DOWNTO 0);
	 SIGNAL  round_bit :	STD_LOGIC;
	 SIGNAL  select_bias_out_2_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  select_bias_out_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  sticky_bits :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  underflow_w :	STD_LOGIC;
	 SIGNAL  underflow_zeros_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  value_add_one_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  value_normal_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  value_zero_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_bias_addition_w_range262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_bias_addition_w_range265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_bias_addition_w_range268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_bias_addition_w_range271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_bias_addition_w_range274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_bias_addition_w_range277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_bias_addition_w_range280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_e1_w_range358w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_e1_w_range368w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range7w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range2w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_not_zero_range260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_not_zero_range263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_not_zero_range266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_not_zero_range269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_not_zero_range272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_not_zero_range275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_not_zero_range278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_remainder_j_w_range362w	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_sticky_bits_range405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_sticky_bits_range409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_sticky_bits_range412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_sticky_bits_range415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_w_quotient_accumulate_w_range385w_range386w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 COMPONENT  altsyncram
	 GENERIC 
	 (
		ADDRESS_ACLR_A	:	STRING := "UNUSED";
		ADDRESS_ACLR_B	:	STRING := "NONE";
		ADDRESS_REG_B	:	STRING := "CLOCK1";
		BYTE_SIZE	:	NATURAL := 8;
		BYTEENA_ACLR_A	:	STRING := "UNUSED";
		BYTEENA_ACLR_B	:	STRING := "NONE";
		BYTEENA_REG_B	:	STRING := "CLOCK1";
		CLOCK_ENABLE_CORE_A	:	STRING := "USE_INPUT_CLKEN";
		CLOCK_ENABLE_CORE_B	:	STRING := "USE_INPUT_CLKEN";
		CLOCK_ENABLE_INPUT_A	:	STRING := "NORMAL";
		CLOCK_ENABLE_INPUT_B	:	STRING := "NORMAL";
		CLOCK_ENABLE_OUTPUT_A	:	STRING := "NORMAL";
		CLOCK_ENABLE_OUTPUT_B	:	STRING := "NORMAL";
		ENABLE_ECC	:	STRING := "FALSE";
		IMPLEMENT_IN_LES	:	STRING := "OFF";
		INDATA_ACLR_A	:	STRING := "UNUSED";
		INDATA_ACLR_B	:	STRING := "NONE";
		INDATA_REG_B	:	STRING := "CLOCK1";
		INIT_FILE	:	STRING := "UNUSED";
		INIT_FILE_LAYOUT	:	STRING := "PORT_A";
		MAXIMUM_DEPTH	:	NATURAL := 0;
		NUMWORDS_A	:	NATURAL := 0;
		NUMWORDS_B	:	NATURAL := 0;
		OPERATION_MODE	:	STRING := "BIDIR_DUAL_PORT";
		OUTDATA_ACLR_A	:	STRING := "NONE";
		OUTDATA_ACLR_B	:	STRING := "NONE";
		OUTDATA_REG_A	:	STRING := "UNREGISTERED";
		OUTDATA_REG_B	:	STRING := "UNREGISTERED";
		POWER_UP_UNINITIALIZED	:	STRING := "FALSE";
		RAM_BLOCK_TYPE	:	STRING := "AUTO";
		RDCONTROL_ACLR_B	:	STRING := "NONE";
		RDCONTROL_REG_B	:	STRING := "CLOCK1";
		READ_DURING_WRITE_MODE_MIXED_PORTS	:	STRING := "DONT_CARE";
		read_during_write_mode_port_a	:	STRING := "NEW_DATA_NO_NBE_READ";
		read_during_write_mode_port_b	:	STRING := "NEW_DATA_NO_NBE_READ";
		WIDTH_A	:	NATURAL;
		WIDTH_B	:	NATURAL := 1;
		WIDTH_BYTEENA_A	:	NATURAL := 1;
		WIDTH_BYTEENA_B	:	NATURAL := 1;
		WIDTH_ECCSTATUS	:	NATURAL := 3;
		WIDTHAD_A	:	NATURAL;
		WIDTHAD_B	:	NATURAL := 1;
		WRCONTROL_ACLR_A	:	STRING := "UNUSED";
		WRCONTROL_ACLR_B	:	STRING := "NONE";
		WRCONTROL_WRADDRESS_REG_B	:	STRING := "CLOCK1";
		INTENDED_DEVICE_FAMILY	:	STRING := "Cyclone II";
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "altsyncram"
	 );
	 PORT
	 ( 
		aclr0	:	IN STD_LOGIC := '0';
		aclr1	:	IN STD_LOGIC := '0';
		address_a	:	IN STD_LOGIC_VECTOR(WIDTHAD_A-1 DOWNTO 0);
		address_b	:	IN STD_LOGIC_VECTOR(WIDTHAD_B-1 DOWNTO 0) := (OTHERS => '1');
		addressstall_a	:	IN STD_LOGIC := '0';
		addressstall_b	:	IN STD_LOGIC := '0';
		byteena_a	:	IN STD_LOGIC_VECTOR(WIDTH_BYTEENA_A-1 DOWNTO 0) := (OTHERS => '1');
		byteena_b	:	IN STD_LOGIC_VECTOR(WIDTH_BYTEENA_B-1 DOWNTO 0) := (OTHERS => '1');
		clock0	:	IN STD_LOGIC := '1';
		clock1	:	IN STD_LOGIC := '1';
		clocken0	:	IN STD_LOGIC := '1';
		clocken1	:	IN STD_LOGIC := '1';
		clocken2	:	IN STD_LOGIC := '1';
		clocken3	:	IN STD_LOGIC := '1';
		data_a	:	IN STD_LOGIC_VECTOR(WIDTH_A-1 DOWNTO 0) := (OTHERS => '1');
		data_b	:	IN STD_LOGIC_VECTOR(WIDTH_B-1 DOWNTO 0) := (OTHERS => '1');
		eccstatus	:	OUT STD_LOGIC_VECTOR(WIDTH_ECCSTATUS-1 DOWNTO 0);
		q_a	:	OUT STD_LOGIC_VECTOR(WIDTH_A-1 DOWNTO 0);
		q_b	:	OUT STD_LOGIC_VECTOR(WIDTH_B-1 DOWNTO 0);
		rden_a	:	IN STD_LOGIC := '1';
		rden_b	:	IN STD_LOGIC := '1';
		wren_a	:	IN STD_LOGIC := '0';
		wren_b	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop0 : FOR i IN 0 TO 7 GENERATE 
		wire_altfp_div_pst1_w_lg_w_lg_w_lg_bias_addition_overf_w304w305w306w(i) <= wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w304w305w(0) AND bias_addition_w(i);
	END GENERATE loop0;
	wire_altfp_div_pst1_w322w(0) <= wire_altfp_div_pst1_w_lg_w_exp_add_output_all_one_range297w321w(0) AND wire_altfp_div_pst1_w_lg_exp_sign_w303w(0);
	wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w304w305w(0) <= wire_altfp_div_pst1_w_lg_bias_addition_overf_w304w(0) AND wire_altfp_div_pst1_w_lg_exp_sign_w303w(0);
	wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w304w312w(0) <= wire_altfp_div_pst1_w_lg_bias_addition_overf_w304w(0) AND exp_sign_w;
	loop1 : FOR i IN 0 TO 7 GENERATE 
		wire_altfp_div_pst1_w302w(i) <= wire_altfp_div_pst1_w_lg_w_lg_w_lg_bias_addition_overf_w299w300w301w(0) AND overflow_ones_w(i);
	END GENERATE loop1;
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range262w286w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range262w(0) AND wire_altfp_div_pst1_w_exp_add_output_all_one_range283w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range265w288w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range265w(0) AND wire_altfp_div_pst1_w_exp_add_output_all_one_range285w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range268w290w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range268w(0) AND wire_altfp_div_pst1_w_exp_add_output_all_one_range287w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range271w292w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range271w(0) AND wire_altfp_div_pst1_w_exp_add_output_all_one_range289w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range274w294w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range274w(0) AND wire_altfp_div_pst1_w_exp_add_output_all_one_range291w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range277w296w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range277w(0) AND wire_altfp_div_pst1_w_exp_add_output_all_one_range293w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range280w298w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range280w(0) AND wire_altfp_div_pst1_w_exp_add_output_all_one_range295w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range11w18w(0) <= wire_altfp_div_pst1_w_dataa_range11w(0) AND wire_altfp_div_pst1_w_exp_a_all_one_w_range7w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range21w28w(0) <= wire_altfp_div_pst1_w_dataa_range21w(0) AND wire_altfp_div_pst1_w_exp_a_all_one_w_range17w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range31w38w(0) <= wire_altfp_div_pst1_w_dataa_range31w(0) AND wire_altfp_div_pst1_w_exp_a_all_one_w_range27w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range41w48w(0) <= wire_altfp_div_pst1_w_dataa_range41w(0) AND wire_altfp_div_pst1_w_exp_a_all_one_w_range37w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range51w58w(0) <= wire_altfp_div_pst1_w_dataa_range51w(0) AND wire_altfp_div_pst1_w_exp_a_all_one_w_range47w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range61w68w(0) <= wire_altfp_div_pst1_w_dataa_range61w(0) AND wire_altfp_div_pst1_w_exp_a_all_one_w_range57w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range71w78w(0) <= wire_altfp_div_pst1_w_dataa_range71w(0) AND wire_altfp_div_pst1_w_exp_a_all_one_w_range67w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range14w20w(0) <= wire_altfp_div_pst1_w_datab_range14w(0) AND wire_altfp_div_pst1_w_exp_b_all_one_w_range9w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range24w30w(0) <= wire_altfp_div_pst1_w_datab_range24w(0) AND wire_altfp_div_pst1_w_exp_b_all_one_w_range19w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range34w40w(0) <= wire_altfp_div_pst1_w_datab_range34w(0) AND wire_altfp_div_pst1_w_exp_b_all_one_w_range29w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range44w50w(0) <= wire_altfp_div_pst1_w_datab_range44w(0) AND wire_altfp_div_pst1_w_exp_b_all_one_w_range39w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range54w60w(0) <= wire_altfp_div_pst1_w_datab_range54w(0) AND wire_altfp_div_pst1_w_exp_b_all_one_w_range49w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range64w70w(0) <= wire_altfp_div_pst1_w_datab_range64w(0) AND wire_altfp_div_pst1_w_exp_b_all_one_w_range59w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range74w80w(0) <= wire_altfp_div_pst1_w_datab_range74w(0) AND wire_altfp_div_pst1_w_exp_b_all_one_w_range69w(0);
	wire_altfp_div_pst1_w_lg_w_exp_a_all_one_w_range77w222w(0) <= wire_altfp_div_pst1_w_exp_a_all_one_w_range77w(0) AND wire_altfp_div_pst1_w_lg_w_man_a_not_zero_w_range214w221w(0);
	wire_altfp_div_pst1_w_lg_w_exp_add_output_all_one_range297w321w(0) <= wire_altfp_div_pst1_w_exp_add_output_all_one_range297w(0) AND wire_altfp_div_pst1_w_lg_bias_addition_overf_w304w(0);
	wire_altfp_div_pst1_w_lg_w_exp_b_all_one_w_range79w224w(0) <= wire_altfp_div_pst1_w_exp_b_all_one_w_range79w(0) AND wire_altfp_div_pst1_w_lg_w_man_b_not_zero_w_range217w223w(0);
	wire_altfp_div_pst1_w_lg_w_exp_b_not_zero_w_range75w256w(0) <= wire_altfp_div_pst1_w_exp_b_not_zero_w_range75w(0) AND wire_altfp_div_pst1_w_lg_w_exp_a_not_zero_w_range72w227w(0);
	wire_altfp_div_pst1_w_lg_a_is_infinity_w233w(0) <= NOT a_is_infinity_w;
	wire_altfp_div_pst1_w_lg_a_is_nan_w234w(0) <= NOT a_is_nan_w;
	wire_altfp_div_pst1_w_lg_bias_addition_overf_w304w(0) <= NOT bias_addition_overf_w;
	wire_altfp_div_pst1_w_lg_exp_sign_w303w(0) <= NOT exp_sign_w;
	wire_altfp_div_pst1_w_lg_w_exp_a_not_zero_w_range72w227w(0) <= NOT wire_altfp_div_pst1_w_exp_a_not_zero_w_range72w(0);
	wire_altfp_div_pst1_w_lg_w_man_a_not_zero_w_range214w221w(0) <= NOT wire_altfp_div_pst1_w_man_a_not_zero_w_range214w(0);
	wire_altfp_div_pst1_w_lg_w_man_b_not_zero_w_range217w223w(0) <= NOT wire_altfp_div_pst1_w_man_b_not_zero_w_range217w(0);
	wire_altfp_div_pst1_w_lg_w_lg_w_lg_bias_addition_overf_w299w300w301w(0) <= wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w299w300w(0) OR a_is_infinity_dffe_1;
	wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w299w300w(0) <= wire_altfp_div_pst1_w_lg_bias_addition_overf_w299w(0) OR nan_pipe_dffe_1;
	wire_altfp_div_pst1_w_lg_bias_addition_overf_w323w(0) <= bias_addition_overf_w OR wire_altfp_div_pst1_w322w(0);
	wire_altfp_div_pst1_w_lg_bias_addition_overf_w299w(0) <= bias_addition_overf_w OR divbyzero_pipe_dffe_1;
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range262w264w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range262w(0) OR wire_altfp_div_pst1_w_exp_add_output_not_zero_range260w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range265w267w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range265w(0) OR wire_altfp_div_pst1_w_exp_add_output_not_zero_range263w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range268w270w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range268w(0) OR wire_altfp_div_pst1_w_exp_add_output_not_zero_range266w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range271w273w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range271w(0) OR wire_altfp_div_pst1_w_exp_add_output_not_zero_range269w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range274w276w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range274w(0) OR wire_altfp_div_pst1_w_exp_add_output_not_zero_range272w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range277w279w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range277w(0) OR wire_altfp_div_pst1_w_exp_add_output_not_zero_range275w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range280w282w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range280w(0) OR wire_altfp_div_pst1_w_exp_add_output_not_zero_range278w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range141w143w(0) <= wire_altfp_div_pst1_w_dataa_range141w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range136w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range147w149w(0) <= wire_altfp_div_pst1_w_dataa_range147w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range142w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range153w155w(0) <= wire_altfp_div_pst1_w_dataa_range153w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range148w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range159w161w(0) <= wire_altfp_div_pst1_w_dataa_range159w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range154w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range165w167w(0) <= wire_altfp_div_pst1_w_dataa_range165w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range160w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range171w173w(0) <= wire_altfp_div_pst1_w_dataa_range171w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range166w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range177w179w(0) <= wire_altfp_div_pst1_w_dataa_range177w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range172w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range183w185w(0) <= wire_altfp_div_pst1_w_dataa_range183w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range178w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range189w191w(0) <= wire_altfp_div_pst1_w_dataa_range189w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range184w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range195w197w(0) <= wire_altfp_div_pst1_w_dataa_range195w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range190w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range87w89w(0) <= wire_altfp_div_pst1_w_dataa_range87w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range82w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range201w203w(0) <= wire_altfp_div_pst1_w_dataa_range201w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range196w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range207w209w(0) <= wire_altfp_div_pst1_w_dataa_range207w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range202w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range213w215w(0) <= wire_altfp_div_pst1_w_dataa_range213w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range208w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range11w13w(0) <= wire_altfp_div_pst1_w_dataa_range11w(0) OR wire_altfp_div_pst1_w_exp_a_not_zero_w_range2w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range21w23w(0) <= wire_altfp_div_pst1_w_dataa_range21w(0) OR wire_altfp_div_pst1_w_exp_a_not_zero_w_range12w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range31w33w(0) <= wire_altfp_div_pst1_w_dataa_range31w(0) OR wire_altfp_div_pst1_w_exp_a_not_zero_w_range22w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range41w43w(0) <= wire_altfp_div_pst1_w_dataa_range41w(0) OR wire_altfp_div_pst1_w_exp_a_not_zero_w_range32w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range51w53w(0) <= wire_altfp_div_pst1_w_dataa_range51w(0) OR wire_altfp_div_pst1_w_exp_a_not_zero_w_range42w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range61w63w(0) <= wire_altfp_div_pst1_w_dataa_range61w(0) OR wire_altfp_div_pst1_w_exp_a_not_zero_w_range52w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range93w95w(0) <= wire_altfp_div_pst1_w_dataa_range93w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range88w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range71w73w(0) <= wire_altfp_div_pst1_w_dataa_range71w(0) OR wire_altfp_div_pst1_w_exp_a_not_zero_w_range62w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range99w101w(0) <= wire_altfp_div_pst1_w_dataa_range99w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range94w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range105w107w(0) <= wire_altfp_div_pst1_w_dataa_range105w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range100w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range111w113w(0) <= wire_altfp_div_pst1_w_dataa_range111w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range106w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range117w119w(0) <= wire_altfp_div_pst1_w_dataa_range117w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range112w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range123w125w(0) <= wire_altfp_div_pst1_w_dataa_range123w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range118w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range129w131w(0) <= wire_altfp_div_pst1_w_dataa_range129w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range124w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range135w137w(0) <= wire_altfp_div_pst1_w_dataa_range135w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range130w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range144w146w(0) <= wire_altfp_div_pst1_w_datab_range144w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range139w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range150w152w(0) <= wire_altfp_div_pst1_w_datab_range150w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range145w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range156w158w(0) <= wire_altfp_div_pst1_w_datab_range156w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range151w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range162w164w(0) <= wire_altfp_div_pst1_w_datab_range162w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range157w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range168w170w(0) <= wire_altfp_div_pst1_w_datab_range168w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range163w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range174w176w(0) <= wire_altfp_div_pst1_w_datab_range174w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range169w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range180w182w(0) <= wire_altfp_div_pst1_w_datab_range180w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range175w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range186w188w(0) <= wire_altfp_div_pst1_w_datab_range186w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range181w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range192w194w(0) <= wire_altfp_div_pst1_w_datab_range192w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range187w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range198w200w(0) <= wire_altfp_div_pst1_w_datab_range198w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range193w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range90w92w(0) <= wire_altfp_div_pst1_w_datab_range90w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range85w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range204w206w(0) <= wire_altfp_div_pst1_w_datab_range204w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range199w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range210w212w(0) <= wire_altfp_div_pst1_w_datab_range210w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range205w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range216w218w(0) <= wire_altfp_div_pst1_w_datab_range216w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range211w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range14w16w(0) <= wire_altfp_div_pst1_w_datab_range14w(0) OR wire_altfp_div_pst1_w_exp_b_not_zero_w_range5w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range24w26w(0) <= wire_altfp_div_pst1_w_datab_range24w(0) OR wire_altfp_div_pst1_w_exp_b_not_zero_w_range15w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range34w36w(0) <= wire_altfp_div_pst1_w_datab_range34w(0) OR wire_altfp_div_pst1_w_exp_b_not_zero_w_range25w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range44w46w(0) <= wire_altfp_div_pst1_w_datab_range44w(0) OR wire_altfp_div_pst1_w_exp_b_not_zero_w_range35w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range54w56w(0) <= wire_altfp_div_pst1_w_datab_range54w(0) OR wire_altfp_div_pst1_w_exp_b_not_zero_w_range45w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range64w66w(0) <= wire_altfp_div_pst1_w_datab_range64w(0) OR wire_altfp_div_pst1_w_exp_b_not_zero_w_range55w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range96w98w(0) <= wire_altfp_div_pst1_w_datab_range96w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range91w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range74w76w(0) <= wire_altfp_div_pst1_w_datab_range74w(0) OR wire_altfp_div_pst1_w_exp_b_not_zero_w_range65w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range102w104w(0) <= wire_altfp_div_pst1_w_datab_range102w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range97w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range108w110w(0) <= wire_altfp_div_pst1_w_datab_range108w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range103w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range114w116w(0) <= wire_altfp_div_pst1_w_datab_range114w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range109w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range120w122w(0) <= wire_altfp_div_pst1_w_datab_range120w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range115w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range126w128w(0) <= wire_altfp_div_pst1_w_datab_range126w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range121w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range132w134w(0) <= wire_altfp_div_pst1_w_datab_range132w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range127w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range138w140w(0) <= wire_altfp_div_pst1_w_datab_range138w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range133w(0);
	a_is_infinity_w <= wire_altfp_div_pst1_w_lg_w_exp_a_all_one_w_range77w222w(0);
	a_is_nan_w <= (exp_a_all_one_w(7) AND man_a_not_zero_w(22));
	a_zero_b_not <= wire_altfp_div_pst1_w_lg_w_exp_b_not_zero_w_range75w256w(0);
	b1_dffe_w <= ( b1_dffe_1);
	b_is_infinity_w <= wire_altfp_div_pst1_w_lg_w_exp_b_all_one_w_range79w224w(0);
	b_is_nan_w <= (exp_b_all_one_w(7) AND man_b_not_zero_w(22));
	bias_addition_overf_w <= wire_bias_addition_overflow;
	bias_addition_w <= wire_bias_addition_result(7 DOWNTO 0);
	both_exp_zeros <= both_exp_zeros_dffe;
	e0_dffe1_wo <= e0_w;
	e0_w <= wire_altsyncram3_q_a;
	e1_w <= ( e1_dffe_1 & e1_dffe_perf_3 & wire_b1_prod_w_lg_w_result_range359w360w);
	exp_a_all_one_w <= ( wire_altfp_div_pst1_w_lg_w_dataa_range71w78w & wire_altfp_div_pst1_w_lg_w_dataa_range61w68w & wire_altfp_div_pst1_w_lg_w_dataa_range51w58w & wire_altfp_div_pst1_w_lg_w_dataa_range41w48w & wire_altfp_div_pst1_w_lg_w_dataa_range31w38w & wire_altfp_div_pst1_w_lg_w_dataa_range21w28w & wire_altfp_div_pst1_w_lg_w_dataa_range11w18w & dataa(23));
	exp_a_not_zero_w <= ( wire_altfp_div_pst1_w_lg_w_dataa_range71w73w & wire_altfp_div_pst1_w_lg_w_dataa_range61w63w & wire_altfp_div_pst1_w_lg_w_dataa_range51w53w & wire_altfp_div_pst1_w_lg_w_dataa_range41w43w & wire_altfp_div_pst1_w_lg_w_dataa_range31w33w & wire_altfp_div_pst1_w_lg_w_dataa_range21w23w & wire_altfp_div_pst1_w_lg_w_dataa_range11w13w & dataa(23));
	exp_add_output_all_one <= ( wire_altfp_div_pst1_w_lg_w_bias_addition_w_range280w298w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range277w296w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range274w294w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range271w292w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range268w290w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range265w288w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range262w286w & bias_addition_w(0));
	exp_add_output_not_zero <= ( wire_altfp_div_pst1_w_lg_w_bias_addition_w_range280w282w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range277w279w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range274w276w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range271w273w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range268w270w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range265w267w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range262w264w & bias_addition_w(0));
	exp_b_all_one_w <= ( wire_altfp_div_pst1_w_lg_w_datab_range74w80w & wire_altfp_div_pst1_w_lg_w_datab_range64w70w & wire_altfp_div_pst1_w_lg_w_datab_range54w60w & wire_altfp_div_pst1_w_lg_w_datab_range44w50w & wire_altfp_div_pst1_w_lg_w_datab_range34w40w & wire_altfp_div_pst1_w_lg_w_datab_range24w30w & wire_altfp_div_pst1_w_lg_w_datab_range14w20w & datab(23));
	exp_b_not_zero_w <= ( wire_altfp_div_pst1_w_lg_w_datab_range74w76w & wire_altfp_div_pst1_w_lg_w_datab_range64w66w & wire_altfp_div_pst1_w_lg_w_datab_range54w56w & wire_altfp_div_pst1_w_lg_w_datab_range44w46w & wire_altfp_div_pst1_w_lg_w_datab_range34w36w & wire_altfp_div_pst1_w_lg_w_datab_range24w26w & wire_altfp_div_pst1_w_lg_w_datab_range14w16w & datab(23));
	exp_result_mux_out <= wire_exp_result_muxa_dataout;
	exp_result_mux_sel_w <= ((((a_zero_b_not_dffe_1 OR b_is_infinity_dffe_1) OR wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w304w312w(0)) OR (((NOT exp_add_output_not_zero(7)) AND wire_altfp_div_pst1_w_lg_bias_addition_overf_w304w(0)) AND wire_altfp_div_pst1_w_lg_exp_sign_w303w(0))) AND wire_nan_pipe_dffe_1_w_lg_q308w(0));
	exp_result_w <= (wire_altfp_div_pst1_w_lg_w_lg_w_lg_bias_addition_overf_w304w305w306w OR wire_altfp_div_pst1_w302w);
	exp_sign_w <= wire_bias_addition_result(8);
	exp_sub_a_w <= ( "0" & dataa(30 DOWNTO 23));
	exp_sub_b_w <= ( "0" & datab(30 DOWNTO 23));
	exp_sub_w <= wire_exp_sub_result;
	frac_a_smaller_dffe1_wi <= frac_a_smaller_w;
	frac_a_smaller_dffe1_wo <= frac_a_smaller_dffe1;
	frac_a_smaller_w <= wire_cmpr2_alb;
	guard_bit <= q_partial_perf_dffe_1(22);
	man_a_adjusted_w <= wire_man_a_adjusteda_dataout;
	man_a_dffe1_wi <= dataa(22 DOWNTO 0);
	man_a_dffe1_wo <= man_a_dffe1_dffe1;
	man_a_not_zero_w <= ( wire_altfp_div_pst1_w_lg_w_dataa_range213w215w & wire_altfp_div_pst1_w_lg_w_dataa_range207w209w & wire_altfp_div_pst1_w_lg_w_dataa_range201w203w & wire_altfp_div_pst1_w_lg_w_dataa_range195w197w & wire_altfp_div_pst1_w_lg_w_dataa_range189w191w & wire_altfp_div_pst1_w_lg_w_dataa_range183w185w & wire_altfp_div_pst1_w_lg_w_dataa_range177w179w & wire_altfp_div_pst1_w_lg_w_dataa_range171w173w & wire_altfp_div_pst1_w_lg_w_dataa_range165w167w & wire_altfp_div_pst1_w_lg_w_dataa_range159w161w & wire_altfp_div_pst1_w_lg_w_dataa_range153w155w & wire_altfp_div_pst1_w_lg_w_dataa_range147w149w & wire_altfp_div_pst1_w_lg_w_dataa_range141w143w & wire_altfp_div_pst1_w_lg_w_dataa_range135w137w & wire_altfp_div_pst1_w_lg_w_dataa_range129w131w & wire_altfp_div_pst1_w_lg_w_dataa_range123w125w & wire_altfp_div_pst1_w_lg_w_dataa_range117w119w & wire_altfp_div_pst1_w_lg_w_dataa_range111w113w & wire_altfp_div_pst1_w_lg_w_dataa_range105w107w & wire_altfp_div_pst1_w_lg_w_dataa_range99w101w & wire_altfp_div_pst1_w_lg_w_dataa_range93w95w & wire_altfp_div_pst1_w_lg_w_dataa_range87w89w & dataa(0));
	man_b_adjusted_w <= ( "1" & man_b_dffe1_wo);
	man_b_dffe1_wi <= datab(22 DOWNTO 0);
	man_b_dffe1_wo <= man_b_dffe1_dffe1;
	man_b_not_zero_w <= ( wire_altfp_div_pst1_w_lg_w_datab_range216w218w & wire_altfp_div_pst1_w_lg_w_datab_range210w212w & wire_altfp_div_pst1_w_lg_w_datab_range204w206w & wire_altfp_div_pst1_w_lg_w_datab_range198w200w & wire_altfp_div_pst1_w_lg_w_datab_range192w194w & wire_altfp_div_pst1_w_lg_w_datab_range186w188w & wire_altfp_div_pst1_w_lg_w_datab_range180w182w & wire_altfp_div_pst1_w_lg_w_datab_range174w176w & wire_altfp_div_pst1_w_lg_w_datab_range168w170w & wire_altfp_div_pst1_w_lg_w_datab_range162w164w & wire_altfp_div_pst1_w_lg_w_datab_range156w158w & wire_altfp_div_pst1_w_lg_w_datab_range150w152w & wire_altfp_div_pst1_w_lg_w_datab_range144w146w & wire_altfp_div_pst1_w_lg_w_datab_range138w140w & wire_altfp_div_pst1_w_lg_w_datab_range132w134w & wire_altfp_div_pst1_w_lg_w_datab_range126w128w & wire_altfp_div_pst1_w_lg_w_datab_range120w122w & wire_altfp_div_pst1_w_lg_w_datab_range114w116w & wire_altfp_div_pst1_w_lg_w_datab_range108w110w & wire_altfp_div_pst1_w_lg_w_datab_range102w104w & wire_altfp_div_pst1_w_lg_w_datab_range96w98w & wire_altfp_div_pst1_w_lg_w_datab_range90w92w & datab(0));
	man_result_dffe_wi <= man_result_w;
	man_result_dffe_wo <= man_result_dffe;
	man_result_mux_select <= (((((over_under_dffe_10 OR a_zero_b_not_dffe_12) OR nan_pipe_dffe_12) OR b_is_infinity_dffe_12) OR a_is_infinity_dffe_12) OR divbyzero_pipe_dffe_12);
	man_result_w <= wire_man_result_muxa_dataout;
	man_zeros_w <= (OTHERS => '0');
	overflow_ones_w <= (OTHERS => '1');
	overflow_underflow <= (overflow_w OR underflow_w);
	overflow_w <= (wire_altfp_div_pst1_w_lg_bias_addition_overf_w323w(0) AND ((wire_nan_pipe_dffe_1_w_lg_q308w(0) AND wire_a_is_infinity_dffe_1_w_lg_q318w(0)) AND wire_divbyzero_pipe_dffe_1_w_lg_q317w(0)));
	quotient_accumulate_w <= ( quotient_k_dffe_0 & "00000000000000" & quotient_j_dffe & "00000000000000");
	quotient_process_cin_w <= (round_bit AND (guard_bit OR sticky_bits(4)));
	remainder_j_w <= ( wire_remainder_sub_0_result(35 DOWNTO 0) & "00000000000000" & wire_a1_prod_result(34 DOWNTO 0) & "000000000000000");
	result <= ( sign_pipe_dffe_13 & exp_result_dffe_11 & man_result_dffe_wo);
	round_bit <= q_partial_perf_dffe_1(21);
	select_bias_out_2_w <= wire_select_bias_2a_dataout;
	select_bias_out_w <= wire_select_biasa_dataout;
	sticky_bits <= ( wire_q_partial_perf_dffe_1_w_lg_w_q_range416w417w & wire_q_partial_perf_dffe_1_w_lg_w_q_range413w414w & wire_q_partial_perf_dffe_1_w_lg_w_q_range410w411w & wire_q_partial_perf_dffe_1_w_lg_w_q_range407w408w & q_partial_perf_dffe_1(16));
	underflow_w <= ((((wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w304w312w(0) OR (((NOT exp_add_output_not_zero(7)) AND wire_altfp_div_pst1_w_lg_bias_addition_overf_w304w(0)) AND wire_altfp_div_pst1_w_lg_exp_sign_w303w(0))) AND wire_nan_pipe_dffe_1_w_lg_q308w(0)) AND wire_a_zero_b_not_dffe_1_w_lg_q326w(0)) AND wire_b_is_infinity_dffe_1_w_lg_q325w(0));
	underflow_zeros_w <= (OTHERS => '0');
	value_add_one_w <= "001111111";
	value_normal_w <= "001111110";
	value_zero_w <= (OTHERS => '0');
	wire_altfp_div_pst1_w_bias_addition_w_range262w(0) <= bias_addition_w(1);
	wire_altfp_div_pst1_w_bias_addition_w_range265w(0) <= bias_addition_w(2);
	wire_altfp_div_pst1_w_bias_addition_w_range268w(0) <= bias_addition_w(3);
	wire_altfp_div_pst1_w_bias_addition_w_range271w(0) <= bias_addition_w(4);
	wire_altfp_div_pst1_w_bias_addition_w_range274w(0) <= bias_addition_w(5);
	wire_altfp_div_pst1_w_bias_addition_w_range277w(0) <= bias_addition_w(6);
	wire_altfp_div_pst1_w_bias_addition_w_range280w(0) <= bias_addition_w(7);
	wire_altfp_div_pst1_w_dataa_range141w(0) <= dataa(10);
	wire_altfp_div_pst1_w_dataa_range147w(0) <= dataa(11);
	wire_altfp_div_pst1_w_dataa_range153w(0) <= dataa(12);
	wire_altfp_div_pst1_w_dataa_range159w(0) <= dataa(13);
	wire_altfp_div_pst1_w_dataa_range165w(0) <= dataa(14);
	wire_altfp_div_pst1_w_dataa_range171w(0) <= dataa(15);
	wire_altfp_div_pst1_w_dataa_range177w(0) <= dataa(16);
	wire_altfp_div_pst1_w_dataa_range183w(0) <= dataa(17);
	wire_altfp_div_pst1_w_dataa_range189w(0) <= dataa(18);
	wire_altfp_div_pst1_w_dataa_range195w(0) <= dataa(19);
	wire_altfp_div_pst1_w_dataa_range87w(0) <= dataa(1);
	wire_altfp_div_pst1_w_dataa_range201w(0) <= dataa(20);
	wire_altfp_div_pst1_w_dataa_range207w(0) <= dataa(21);
	wire_altfp_div_pst1_w_dataa_range213w(0) <= dataa(22);
	wire_altfp_div_pst1_w_dataa_range11w(0) <= dataa(24);
	wire_altfp_div_pst1_w_dataa_range21w(0) <= dataa(25);
	wire_altfp_div_pst1_w_dataa_range31w(0) <= dataa(26);
	wire_altfp_div_pst1_w_dataa_range41w(0) <= dataa(27);
	wire_altfp_div_pst1_w_dataa_range51w(0) <= dataa(28);
	wire_altfp_div_pst1_w_dataa_range61w(0) <= dataa(29);
	wire_altfp_div_pst1_w_dataa_range93w(0) <= dataa(2);
	wire_altfp_div_pst1_w_dataa_range71w(0) <= dataa(30);
	wire_altfp_div_pst1_w_dataa_range99w(0) <= dataa(3);
	wire_altfp_div_pst1_w_dataa_range105w(0) <= dataa(4);
	wire_altfp_div_pst1_w_dataa_range111w(0) <= dataa(5);
	wire_altfp_div_pst1_w_dataa_range117w(0) <= dataa(6);
	wire_altfp_div_pst1_w_dataa_range123w(0) <= dataa(7);
	wire_altfp_div_pst1_w_dataa_range129w(0) <= dataa(8);
	wire_altfp_div_pst1_w_dataa_range135w(0) <= dataa(9);
	wire_altfp_div_pst1_w_datab_range144w(0) <= datab(10);
	wire_altfp_div_pst1_w_datab_range150w(0) <= datab(11);
	wire_altfp_div_pst1_w_datab_range156w(0) <= datab(12);
	wire_altfp_div_pst1_w_datab_range162w(0) <= datab(13);
	wire_altfp_div_pst1_w_datab_range168w(0) <= datab(14);
	wire_altfp_div_pst1_w_datab_range174w(0) <= datab(15);
	wire_altfp_div_pst1_w_datab_range180w(0) <= datab(16);
	wire_altfp_div_pst1_w_datab_range186w(0) <= datab(17);
	wire_altfp_div_pst1_w_datab_range192w(0) <= datab(18);
	wire_altfp_div_pst1_w_datab_range198w(0) <= datab(19);
	wire_altfp_div_pst1_w_datab_range90w(0) <= datab(1);
	wire_altfp_div_pst1_w_datab_range204w(0) <= datab(20);
	wire_altfp_div_pst1_w_datab_range210w(0) <= datab(21);
	wire_altfp_div_pst1_w_datab_range216w(0) <= datab(22);
	wire_altfp_div_pst1_w_datab_range14w(0) <= datab(24);
	wire_altfp_div_pst1_w_datab_range24w(0) <= datab(25);
	wire_altfp_div_pst1_w_datab_range34w(0) <= datab(26);
	wire_altfp_div_pst1_w_datab_range44w(0) <= datab(27);
	wire_altfp_div_pst1_w_datab_range54w(0) <= datab(28);
	wire_altfp_div_pst1_w_datab_range64w(0) <= datab(29);
	wire_altfp_div_pst1_w_datab_range96w(0) <= datab(2);
	wire_altfp_div_pst1_w_datab_range74w(0) <= datab(30);
	wire_altfp_div_pst1_w_datab_range102w(0) <= datab(3);
	wire_altfp_div_pst1_w_datab_range108w(0) <= datab(4);
	wire_altfp_div_pst1_w_datab_range114w(0) <= datab(5);
	wire_altfp_div_pst1_w_datab_range120w(0) <= datab(6);
	wire_altfp_div_pst1_w_datab_range126w(0) <= datab(7);
	wire_altfp_div_pst1_w_datab_range132w(0) <= datab(8);
	wire_altfp_div_pst1_w_datab_range138w(0) <= datab(9);
	wire_altfp_div_pst1_w_e1_w_range358w <= e1_w(16 DOWNTO 0);
	wire_altfp_div_pst1_w_e1_w_range368w <= e1_w(33 DOWNTO 17);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range7w(0) <= exp_a_all_one_w(0);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range17w(0) <= exp_a_all_one_w(1);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range27w(0) <= exp_a_all_one_w(2);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range37w(0) <= exp_a_all_one_w(3);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range47w(0) <= exp_a_all_one_w(4);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range57w(0) <= exp_a_all_one_w(5);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range67w(0) <= exp_a_all_one_w(6);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range77w(0) <= exp_a_all_one_w(7);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range2w(0) <= exp_a_not_zero_w(0);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range12w(0) <= exp_a_not_zero_w(1);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range22w(0) <= exp_a_not_zero_w(2);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range32w(0) <= exp_a_not_zero_w(3);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range42w(0) <= exp_a_not_zero_w(4);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range52w(0) <= exp_a_not_zero_w(5);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range62w(0) <= exp_a_not_zero_w(6);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range72w(0) <= exp_a_not_zero_w(7);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range283w(0) <= exp_add_output_all_one(0);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range285w(0) <= exp_add_output_all_one(1);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range287w(0) <= exp_add_output_all_one(2);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range289w(0) <= exp_add_output_all_one(3);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range291w(0) <= exp_add_output_all_one(4);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range293w(0) <= exp_add_output_all_one(5);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range295w(0) <= exp_add_output_all_one(6);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range297w(0) <= exp_add_output_all_one(7);
	wire_altfp_div_pst1_w_exp_add_output_not_zero_range260w(0) <= exp_add_output_not_zero(0);
	wire_altfp_div_pst1_w_exp_add_output_not_zero_range263w(0) <= exp_add_output_not_zero(1);
	wire_altfp_div_pst1_w_exp_add_output_not_zero_range266w(0) <= exp_add_output_not_zero(2);
	wire_altfp_div_pst1_w_exp_add_output_not_zero_range269w(0) <= exp_add_output_not_zero(3);
	wire_altfp_div_pst1_w_exp_add_output_not_zero_range272w(0) <= exp_add_output_not_zero(4);
	wire_altfp_div_pst1_w_exp_add_output_not_zero_range275w(0) <= exp_add_output_not_zero(5);
	wire_altfp_div_pst1_w_exp_add_output_not_zero_range278w(0) <= exp_add_output_not_zero(6);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range9w(0) <= exp_b_all_one_w(0);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range19w(0) <= exp_b_all_one_w(1);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range29w(0) <= exp_b_all_one_w(2);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range39w(0) <= exp_b_all_one_w(3);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range49w(0) <= exp_b_all_one_w(4);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range59w(0) <= exp_b_all_one_w(5);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range69w(0) <= exp_b_all_one_w(6);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range79w(0) <= exp_b_all_one_w(7);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range5w(0) <= exp_b_not_zero_w(0);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range15w(0) <= exp_b_not_zero_w(1);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range25w(0) <= exp_b_not_zero_w(2);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range35w(0) <= exp_b_not_zero_w(3);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range45w(0) <= exp_b_not_zero_w(4);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range55w(0) <= exp_b_not_zero_w(5);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range65w(0) <= exp_b_not_zero_w(6);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range75w(0) <= exp_b_not_zero_w(7);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range82w(0) <= man_a_not_zero_w(0);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range142w(0) <= man_a_not_zero_w(10);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range148w(0) <= man_a_not_zero_w(11);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range154w(0) <= man_a_not_zero_w(12);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range160w(0) <= man_a_not_zero_w(13);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range166w(0) <= man_a_not_zero_w(14);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range172w(0) <= man_a_not_zero_w(15);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range178w(0) <= man_a_not_zero_w(16);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range184w(0) <= man_a_not_zero_w(17);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range190w(0) <= man_a_not_zero_w(18);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range196w(0) <= man_a_not_zero_w(19);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range88w(0) <= man_a_not_zero_w(1);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range202w(0) <= man_a_not_zero_w(20);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range208w(0) <= man_a_not_zero_w(21);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range214w(0) <= man_a_not_zero_w(22);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range94w(0) <= man_a_not_zero_w(2);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range100w(0) <= man_a_not_zero_w(3);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range106w(0) <= man_a_not_zero_w(4);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range112w(0) <= man_a_not_zero_w(5);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range118w(0) <= man_a_not_zero_w(6);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range124w(0) <= man_a_not_zero_w(7);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range130w(0) <= man_a_not_zero_w(8);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range136w(0) <= man_a_not_zero_w(9);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range85w(0) <= man_b_not_zero_w(0);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range145w(0) <= man_b_not_zero_w(10);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range151w(0) <= man_b_not_zero_w(11);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range157w(0) <= man_b_not_zero_w(12);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range163w(0) <= man_b_not_zero_w(13);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range169w(0) <= man_b_not_zero_w(14);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range175w(0) <= man_b_not_zero_w(15);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range181w(0) <= man_b_not_zero_w(16);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range187w(0) <= man_b_not_zero_w(17);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range193w(0) <= man_b_not_zero_w(18);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range199w(0) <= man_b_not_zero_w(19);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range91w(0) <= man_b_not_zero_w(1);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range205w(0) <= man_b_not_zero_w(20);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range211w(0) <= man_b_not_zero_w(21);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range217w(0) <= man_b_not_zero_w(22);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range97w(0) <= man_b_not_zero_w(2);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range103w(0) <= man_b_not_zero_w(3);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range109w(0) <= man_b_not_zero_w(4);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range115w(0) <= man_b_not_zero_w(5);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range121w(0) <= man_b_not_zero_w(6);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range127w(0) <= man_b_not_zero_w(7);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range133w(0) <= man_b_not_zero_w(8);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range139w(0) <= man_b_not_zero_w(9);
	wire_altfp_div_pst1_w_remainder_j_w_range362w <= remainder_j_w(49 DOWNTO 0);
	wire_altfp_div_pst1_w_sticky_bits_range405w(0) <= sticky_bits(0);
	wire_altfp_div_pst1_w_sticky_bits_range409w(0) <= sticky_bits(1);
	wire_altfp_div_pst1_w_sticky_bits_range412w(0) <= sticky_bits(2);
	wire_altfp_div_pst1_w_sticky_bits_range415w(0) <= sticky_bits(3);
	wire_altfp_div_pst1_w_w_quotient_accumulate_w_range385w_range386w <= quotient_accumulate_w(30 DOWNTO 14);
	altsyncram3 :  altsyncram
	  GENERIC MAP (
		INIT_FILE => "k_ukf_div.hex",
		OPERATION_MODE => "ROM",
		WIDTH_A => 9,
		WIDTHAD_A => 9,
		INTENDED_DEVICE_FAMILY => "Cyclone II"
	  )
	  PORT MAP ( 
		address_a => datab(22 DOWNTO 14),
		clock0 => clock,
		clocken0 => clk_en,
		q_a => wire_altsyncram3_q_a
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_0 <= a_is_infinity_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_1 <= a_is_infinity_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	wire_a_is_infinity_dffe_1_w_lg_q318w(0) <= NOT a_is_infinity_dffe_1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_10 <= a_is_infinity_dffe_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_11 <= a_is_infinity_dffe_10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_12 <= a_is_infinity_dffe_11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_2 <= a_is_infinity_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_3 <= a_is_infinity_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_4 <= a_is_infinity_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_5 <= a_is_infinity_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_6 <= a_is_infinity_dffe_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_7 <= a_is_infinity_dffe_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_8 <= a_is_infinity_dffe_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_9 <= a_is_infinity_dffe_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_0 <= a_zero_b_not;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_1 <= a_zero_b_not_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	wire_a_zero_b_not_dffe_1_w_lg_q326w(0) <= NOT a_zero_b_not_dffe_1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_10 <= a_zero_b_not_dffe_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_11 <= a_zero_b_not_dffe_10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_12 <= a_zero_b_not_dffe_11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_2 <= a_zero_b_not_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_3 <= a_zero_b_not_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_4 <= a_zero_b_not_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_5 <= a_zero_b_not_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_6 <= a_zero_b_not_dffe_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_7 <= a_zero_b_not_dffe_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_8 <= a_zero_b_not_dffe_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_9 <= a_zero_b_not_dffe_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b1_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b1_dffe_0 <= wire_b1_prod_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b1_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b1_dffe_1 <= b1_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_0 <= b_is_infinity_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_1 <= b_is_infinity_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	wire_b_is_infinity_dffe_1_w_lg_q325w(0) <= NOT b_is_infinity_dffe_1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_10 <= b_is_infinity_dffe_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_11 <= b_is_infinity_dffe_10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_12 <= b_is_infinity_dffe_11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_2 <= b_is_infinity_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_3 <= b_is_infinity_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_4 <= b_is_infinity_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_5 <= b_is_infinity_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_6 <= b_is_infinity_dffe_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_7 <= b_is_infinity_dffe_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_8 <= b_is_infinity_dffe_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_9 <= b_is_infinity_dffe_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN both_exp_zeros_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN both_exp_zeros_dffe <= ((NOT exp_b_not_zero_w(7)) AND wire_altfp_div_pst1_w_lg_w_exp_a_not_zero_w_range72w227w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_0 <= ((((NOT exp_b_not_zero_w(7)) AND wire_altfp_div_pst1_w_lg_a_is_nan_w234w(0)) AND exp_a_not_zero_w(7)) AND wire_altfp_div_pst1_w_lg_a_is_infinity_w233w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_1 <= divbyzero_pipe_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	wire_divbyzero_pipe_dffe_1_w_lg_q317w(0) <= NOT divbyzero_pipe_dffe_1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_10 <= divbyzero_pipe_dffe_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_11 <= divbyzero_pipe_dffe_10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_12 <= divbyzero_pipe_dffe_11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_2 <= divbyzero_pipe_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_3 <= divbyzero_pipe_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_4 <= divbyzero_pipe_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_5 <= divbyzero_pipe_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_6 <= divbyzero_pipe_dffe_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_7 <= divbyzero_pipe_dffe_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_8 <= divbyzero_pipe_dffe_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_9 <= divbyzero_pipe_dffe_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN e1_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN e1_dffe_0 <= wire_altfp_div_pst1_w_e1_w_range358w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN e1_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN e1_dffe_1 <= wire_altfp_div_pst1_w_e1_w_range368w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN e1_dffe_perf_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN e1_dffe_perf_0 <= e1_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN e1_dffe_perf_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN e1_dffe_perf_1 <= e1_dffe_perf_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN e1_dffe_perf_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN e1_dffe_perf_2 <= e1_dffe_perf_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN e1_dffe_perf_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN e1_dffe_perf_3 <= e1_dffe_perf_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_0 <= exp_result_mux_out;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_1 <= exp_result_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_10 <= exp_result_dffe_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_11 <= exp_result_dffe_10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_2 <= exp_result_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_3 <= exp_result_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_4 <= exp_result_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_5 <= exp_result_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_6 <= exp_result_dffe_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_7 <= exp_result_dffe_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_8 <= exp_result_dffe_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_9 <= exp_result_dffe_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN frac_a_smaller_dffe1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN frac_a_smaller_dffe1 <= frac_a_smaller_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_a_dffe1_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_a_dffe1_dffe1 <= man_a_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_b_dffe1_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_b_dffe1_dffe1 <= man_b_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_result_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_result_dffe <= man_result_dffe_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_0 <= (((a_is_nan_w OR b_is_nan_w) OR (a_is_infinity_w AND b_is_infinity_w)) OR (wire_altfp_div_pst1_w_lg_w_exp_a_not_zero_w_range72w227w(0) AND (NOT exp_b_not_zero_w(7))));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_1 <= nan_pipe_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	wire_nan_pipe_dffe_1_w_lg_q308w(0) <= NOT nan_pipe_dffe_1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_10 <= nan_pipe_dffe_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_11 <= nan_pipe_dffe_10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_12 <= nan_pipe_dffe_11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_2 <= nan_pipe_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_3 <= nan_pipe_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_4 <= nan_pipe_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_5 <= nan_pipe_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_6 <= nan_pipe_dffe_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_7 <= nan_pipe_dffe_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_8 <= nan_pipe_dffe_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_9 <= nan_pipe_dffe_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN over_under_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN over_under_dffe_0 <= overflow_underflow;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN over_under_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN over_under_dffe_1 <= over_under_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN over_under_dffe_10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN over_under_dffe_10 <= over_under_dffe_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN over_under_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN over_under_dffe_2 <= over_under_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN over_under_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN over_under_dffe_3 <= over_under_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN over_under_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN over_under_dffe_4 <= over_under_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN over_under_dffe_5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN over_under_dffe_5 <= over_under_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN over_under_dffe_6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN over_under_dffe_6 <= over_under_dffe_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN over_under_dffe_7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN over_under_dffe_7 <= over_under_dffe_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN over_under_dffe_8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN over_under_dffe_8 <= over_under_dffe_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN over_under_dffe_9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN over_under_dffe_9 <= over_under_dffe_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_partial_perf_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN q_partial_perf_dffe_0 <= wire_q_partial_0_result;
			END IF;
		END IF;
	END PROCESS;
	wire_q_partial_perf_dffe_0_w_q_range373w <= q_partial_perf_dffe_0(32 DOWNTO 16);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_partial_perf_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN q_partial_perf_dffe_1 <= wire_q_partial_1_result;
			END IF;
		END IF;
	END PROCESS;
	wire_q_partial_perf_dffe_1_w_lg_w_q_range407w408w(0) <= wire_q_partial_perf_dffe_1_w_q_range407w(0) OR wire_altfp_div_pst1_w_sticky_bits_range405w(0);
	wire_q_partial_perf_dffe_1_w_lg_w_q_range410w411w(0) <= wire_q_partial_perf_dffe_1_w_q_range410w(0) OR wire_altfp_div_pst1_w_sticky_bits_range409w(0);
	wire_q_partial_perf_dffe_1_w_lg_w_q_range413w414w(0) <= wire_q_partial_perf_dffe_1_w_q_range413w(0) OR wire_altfp_div_pst1_w_sticky_bits_range412w(0);
	wire_q_partial_perf_dffe_1_w_lg_w_q_range416w417w(0) <= wire_q_partial_perf_dffe_1_w_q_range416w(0) OR wire_altfp_div_pst1_w_sticky_bits_range415w(0);
	wire_q_partial_perf_dffe_1_w_q_range407w(0) <= q_partial_perf_dffe_1(17);
	wire_q_partial_perf_dffe_1_w_q_range410w(0) <= q_partial_perf_dffe_1(18);
	wire_q_partial_perf_dffe_1_w_q_range413w(0) <= q_partial_perf_dffe_1(19);
	wire_q_partial_perf_dffe_1_w_q_range416w(0) <= q_partial_perf_dffe_1(20);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN quotient_j_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN quotient_j_dffe <= wire_q_partial_perf_dffe_0_w_q_range373w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN quotient_k_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN quotient_k_dffe_0 <= quotient_k_dffe_perf_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN quotient_k_dffe_perf_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN quotient_k_dffe_perf_0 <= wire_altfp_div_pst1_w_w_quotient_accumulate_w_range385w_range386w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN quotient_k_dffe_perf_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN quotient_k_dffe_perf_1 <= quotient_k_dffe_perf_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN quotient_k_dffe_perf_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN quotient_k_dffe_perf_2 <= quotient_k_dffe_perf_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN quotient_k_dffe_perf_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN quotient_k_dffe_perf_3 <= quotient_k_dffe_perf_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN remainder_j_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN remainder_j_dffe_0 <= wire_altfp_div_pst1_w_remainder_j_w_range362w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN remainder_j_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN remainder_j_dffe_1 <= remainder_j_dffe_perf_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN remainder_j_dffe_perf_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN remainder_j_dffe_perf_0 <= remainder_j_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN remainder_j_dffe_perf_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN remainder_j_dffe_perf_1 <= remainder_j_dffe_perf_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN remainder_j_dffe_perf_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN remainder_j_dffe_perf_2 <= remainder_j_dffe_perf_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_0 <= (dataa(31) XOR datab(31));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_1 <= sign_pipe_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_10 <= sign_pipe_dffe_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_11 <= sign_pipe_dffe_10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_12 <= sign_pipe_dffe_11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_13 <= sign_pipe_dffe_12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_2 <= sign_pipe_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_3 <= sign_pipe_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_4 <= sign_pipe_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_5 <= sign_pipe_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_6 <= sign_pipe_dffe_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_7 <= sign_pipe_dffe_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_8 <= sign_pipe_dffe_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_9 <= sign_pipe_dffe_8;
			END IF;
		END IF;
	END PROCESS;
	bias_addition :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => exp_sub_w,
		datab => select_bias_out_2_w,
		overflow => wire_bias_addition_overflow,
		result => wire_bias_addition_result
	  );
	exp_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => exp_sub_a_w,
		datab => exp_sub_b_w,
		result => wire_exp_sub_result
	  );
	wire_quotient_process_dataa <= ( quotient_accumulate_w(61 DOWNTO 45) & "00000000000000");
	wire_quotient_process_datab <= ( "00000000000000" & q_partial_perf_dffe_1(32 DOWNTO 22) & "111111");
	wire_quotient_process_w_result_range425w <= wire_quotient_process_result(28 DOWNTO 6);
	quotient_process :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 31
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => quotient_process_cin_w,
		clken => clk_en,
		clock => clock,
		dataa => wire_quotient_process_dataa,
		datab => wire_quotient_process_datab,
		result => wire_quotient_process_result
	  );
	wire_remainder_sub_0_dataa <= ( remainder_j_dffe_1(49 DOWNTO 15) & "000000000000000");
	remainder_sub_0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 50
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_remainder_sub_0_dataa,
		datab => wire_remainder_mult_0_result(49 DOWNTO 0),
		result => wire_remainder_sub_0_result
	  );
	cmpr2 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 23
	  )
	  PORT MAP ( 
		alb => wire_cmpr2_alb,
		dataa => dataa(22 DOWNTO 0),
		datab => datab(22 DOWNTO 0)
	  );
	wire_a1_prod_datab <= ( "1" & e0_dffe1_wo);
	a1_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 25,
		LPM_WIDTHB => 10,
		LPM_WIDTHP => 35,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => man_a_adjusted_w,
		datab => wire_a1_prod_datab,
		result => wire_a1_prod_result
	  );
	loop2 : FOR i IN 0 TO 16 GENERATE 
		wire_b1_prod_w_lg_w_result_range359w360w(i) <= NOT wire_b1_prod_w_result_range359w(i);
	END GENERATE loop2;
	wire_b1_prod_datab <= ( "1" & e0_dffe1_wo);
	wire_b1_prod_w_result_range359w <= wire_b1_prod_result(33 DOWNTO 17);
	b1_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 24,
		LPM_WIDTHB => 10,
		LPM_WIDTHP => 34,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => man_b_adjusted_w,
		datab => wire_b1_prod_datab,
		result => wire_b1_prod_result
	  );
	q_partial_0 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 17,
		LPM_WIDTHB => 17,
		LPM_WIDTHP => 34,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => remainder_j_w(49 DOWNTO 33),
		datab => e1_w(16 DOWNTO 0),
		result => wire_q_partial_0_result
	  );
	q_partial_1 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 17,
		LPM_WIDTHB => 17,
		LPM_WIDTHP => 34,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => remainder_j_w(99 DOWNTO 83),
		datab => e1_w(50 DOWNTO 34),
		result => wire_q_partial_1_result
	  );
	remainder_mult_0 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 34,
		LPM_WIDTHB => 17,
		LPM_WIDTHP => 51,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => b1_dffe_w(33 DOWNTO 0),
		datab => q_partial_perf_dffe_0(32 DOWNTO 16),
		result => wire_remainder_mult_0_result
	  );
	wire_exp_result_muxa_dataout <= underflow_zeros_w WHEN exp_result_mux_sel_w = '1'  ELSE exp_result_w;
	wire_man_a_adjusteda_dataout <= ( "1" & man_a_dffe1_wo & "0") WHEN frac_a_smaller_dffe1_wo = '1'  ELSE ( "0" & "1" & man_a_dffe1_wo);
	wire_man_result_muxa_dataout <= ( nan_pipe_dffe_12 & man_zeros_w(21 DOWNTO 0)) WHEN man_result_mux_select = '1'  ELSE wire_quotient_process_result(28 DOWNTO 6);
	wire_select_bias_2a_dataout <= value_zero_w WHEN both_exp_zeros = '1'  ELSE select_bias_out_w;
	wire_select_biasa_dataout <= value_normal_w WHEN frac_a_smaller_dffe1_wo = '1'  ELSE value_add_one_w;

 END RTL; --k_ukf_div_altfp_div_pst_o3f

--synthesis_resources = altsyncram 1 lpm_add_sub 4 lpm_compare 1 lpm_mult 5 mux21 74 reg 847 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  k_ukf_div_altfp_div_79h IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 datab	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END k_ukf_div_altfp_div_79h;

 ARCHITECTURE RTL OF k_ukf_div_altfp_div_79h IS

	 SIGNAL  wire_altfp_div_pst1_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  clk_en	:	STD_LOGIC;
	 COMPONENT  k_ukf_div_altfp_div_pst_o3f
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC;
		dataa	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		datab	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	aclr <= '0';
	clk_en <= '1';
	result <= wire_altfp_div_pst1_result;
	altfp_div_pst1 :  k_ukf_div_altfp_div_pst_o3f
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		dataa => dataa,
		datab => datab,
		result => wire_altfp_div_pst1_result
	  );

 END RTL; --k_ukf_div_altfp_div_79h
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY k_ukf_div IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END k_ukf_div;


ARCHITECTURE RTL OF k_ukf_div IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT k_ukf_div_altfp_div_79h
	PORT (
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	k_ukf_div_altfp_div_79h_component : k_ukf_div_altfp_div_79h
	PORT MAP (
		clock => clock,
		dataa => dataa,
		datab => datab,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "1"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: DENORMAL_SUPPORT STRING "NO"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: CONSTANT: OPTIMIZE STRING "SPEED"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "14"
-- Retrieval info: CONSTANT: REDUCED_FUNCTIONALITY STRING "NO"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: dataa 0 0 32 0 INPUT NODEFVAL "dataa[31..0]"
-- Retrieval info: USED_PORT: datab 0 0 32 0 INPUT NODEFVAL "datab[31..0]"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @dataa 0 0 32 0 dataa 0 0 32 0
-- Retrieval info: CONNECT: @datab 0 0 32 0 datab 0 0 32 0
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL k_ukf_div.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL k_ukf_div.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL k_ukf_div.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL k_ukf_div.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL k_ukf_div_inst.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL k_ukf_div_syn.v TRUE
