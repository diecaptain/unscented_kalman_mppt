-- megafunction wizard: %ALTFP_SQRT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altfp_sqrt 

-- ============================================================
-- File Name: k_ukf_sqrt.vhd
-- Megafunction Name(s):
-- 			altfp_sqrt
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.1 Build 259 01/25/2012 SP 2 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altfp_sqrt CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" PIPELINE=28 ROUNDING="TO_NEAREST" WIDTH_EXP=8 WIDTH_MAN=23 clock data result
--VERSION_BEGIN 11.1SP2 cbx_altfp_sqrt 2012:01:25:21:13:53:SJ cbx_cycloneii 2012:01:25:21:13:53:SJ cbx_lpm_add_sub 2012:01:25:21:13:53:SJ cbx_mgl 2012:01:25:21:15:41:SJ cbx_stratix 2012:01:25:21:13:53:SJ cbx_stratixii 2012:01:25:21:13:53:SJ  VERSION_END


--alt_sqrt_block CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" PIPELINE=28 WIDTH_SQRT=25 aclr clken clock rad root_result
--VERSION_BEGIN 11.1SP2 cbx_altfp_sqrt 2012:01:25:21:13:53:SJ cbx_cycloneii 2012:01:25:21:13:53:SJ cbx_lpm_add_sub 2012:01:25:21:13:53:SJ cbx_mgl 2012:01:25:21:15:41:SJ cbx_stratix 2012:01:25:21:13:53:SJ cbx_stratixii 2012:01:25:21:13:53:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 25 reg 1034 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  k_ukf_sqrt_alt_sqrt_block_nfb IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 rad	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0);
		 root_result	:	OUT  STD_LOGIC_VECTOR (24 DOWNTO 0)
	 ); 
 END k_ukf_sqrt_alt_sqrt_block_nfb;

 ARCHITECTURE RTL OF k_ukf_sqrt_alt_sqrt_block_nfb IS

	 SIGNAL	 q_ff0c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff10c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff11c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff12c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff13c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff14c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff15c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff16c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff17c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff18c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff19c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff1c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff20c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff21c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff22c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff23c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff2c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff3c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff4c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff5c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff6c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff7c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff8c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff9c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rad_ff0c	:	STD_LOGIC_VECTOR(25 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rad_ff10c	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff10c_w_lg_w_lg_w_q_range2589w2592w2593w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_rad_ff10c_w_lg_w_q_range2589w2590w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_rad_ff10c_w_lg_w_q_range2589w2592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff10c_w_lg_w_lg_w_lg_w_q_range2589w2592w2593w2594w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_rad_ff10c_w_q_range2589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff11c	:	STD_LOGIC_VECTOR(14 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff11c_w_lg_w_lg_w_q_range2620w2623w2624w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_rad_ff11c_w_lg_w_q_range2620w2621w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_rad_ff11c_w_lg_w_q_range2620w2623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff11c_w_lg_w_lg_w_lg_w_q_range2620w2623w2624w2625w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_rad_ff11c_w_q_range2620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff12c	:	STD_LOGIC_VECTOR(13 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff12c_w_lg_w_lg_w_q_range2652w2655w2656w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_rad_ff12c_w_lg_w_q_range2652w2653w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_rad_ff12c_w_lg_w_q_range2652w2655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff12c_w_lg_w_lg_w_lg_w_q_range2652w2655w2656w2657w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_rad_ff12c_w_q_range2652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff13c	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff13c_w_lg_w_lg_w_q_range2691w2694w2695w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_rad_ff13c_w_lg_w_q_range2691w2692w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_rad_ff13c_w_lg_w_q_range2691w2694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff13c_w_lg_w_lg_w_lg_w_q_range2691w2694w2695w2696w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_rad_ff13c_w_q_range2691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff14c	:	STD_LOGIC_VECTOR(13 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff14c_w_lg_w_lg_w_q_range2730w2733w2734w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_rad_ff14c_w_lg_w_q_range2730w2731w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_rad_ff14c_w_lg_w_q_range2730w2733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff14c_w_lg_w_lg_w_lg_w_q_range2730w2733w2734w2735w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_rad_ff14c_w_q_range2730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff15c	:	STD_LOGIC_VECTOR(14 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff15c_w_lg_w_lg_w_q_range2769w2772w2773w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_rad_ff15c_w_lg_w_q_range2769w2770w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_rad_ff15c_w_lg_w_q_range2769w2772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff15c_w_lg_w_lg_w_lg_w_q_range2769w2772w2773w2774w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_rad_ff15c_w_q_range2769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff16c	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff16c_w_lg_w_lg_w_q_range2808w2811w2812w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_rad_ff16c_w_lg_w_q_range2808w2809w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_rad_ff16c_w_lg_w_q_range2808w2811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff16c_w_lg_w_lg_w_lg_w_q_range2808w2811w2812w2813w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_rad_ff16c_w_q_range2808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff17c	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff17c_w_lg_w_lg_w_q_range2847w2850w2851w	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_rad_ff17c_w_lg_w_q_range2847w2848w	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_rad_ff17c_w_lg_w_q_range2847w2850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff17c_w_lg_w_lg_w_lg_w_q_range2847w2850w2851w2852w	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_rad_ff17c_w_q_range2847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff18c	:	STD_LOGIC_VECTOR(17 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff18c_w_lg_w_lg_w_q_range2886w2889w2890w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_rad_ff18c_w_lg_w_q_range2886w2887w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_rad_ff18c_w_lg_w_q_range2886w2889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff18c_w_lg_w_lg_w_lg_w_q_range2886w2889w2890w2891w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_rad_ff18c_w_q_range2886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff19c	:	STD_LOGIC_VECTOR(18 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff19c_w_lg_w_lg_w_q_range2925w2928w2929w	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_rad_ff19c_w_lg_w_q_range2925w2926w	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_rad_ff19c_w_lg_w_q_range2925w2928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff19c_w_lg_w_lg_w_lg_w_q_range2925w2928w2929w2930w	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_rad_ff19c_w_q_range2925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff1c	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff1c_w_lg_w_lg_w_q_range2301w2304w2305w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_rad_ff1c_w_lg_w_q_range2301w2302w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_rad_ff1c_w_lg_w_q_range2301w2304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff1c_w_lg_w_lg_w_lg_w_q_range2301w2304w2305w2306w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_rad_ff1c_w_q_range2301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff20c	:	STD_LOGIC_VECTOR(19 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff20c_w_lg_w_lg_w_q_range2964w2967w2968w	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_rad_ff20c_w_lg_w_q_range2964w2965w	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_rad_ff20c_w_lg_w_q_range2964w2967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff20c_w_lg_w_lg_w_lg_w_q_range2964w2967w2968w2969w	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_rad_ff20c_w_q_range2964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff21c	:	STD_LOGIC_VECTOR(20 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff21c_w_lg_w_lg_w_q_range3003w3006w3007w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_rad_ff21c_w_lg_w_q_range3003w3004w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_rad_ff21c_w_lg_w_q_range3003w3006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff21c_w_lg_w_lg_w_lg_w_q_range3003w3006w3007w3008w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_rad_ff21c_w_q_range3003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff22c	:	STD_LOGIC_VECTOR(21 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff22c_w_lg_w_lg_w_q_range3042w3045w3046w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_rad_ff22c_w_lg_w_q_range3042w3043w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_rad_ff22c_w_lg_w_q_range3042w3045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff22c_w_lg_w_lg_w_lg_w_q_range3042w3045w3046w3047w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_rad_ff22c_w_q_range3042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff23c	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff23c_w_lg_w_lg_w_q_range3069w3070w3086w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_rad_ff23c_w_lg_w_q_range3069w3084w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_rad_ff23c_w_lg_w_q_range3069w3070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff23c_w_lg_w_lg_w_lg_w_q_range3069w3070w3086w3087w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_rad_ff23c_w_q_range3069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff2c	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff2c_w_lg_w_lg_w_q_range2333w2336w2337w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_rad_ff2c_w_lg_w_q_range2333w2334w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_rad_ff2c_w_lg_w_q_range2333w2336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff2c_w_lg_w_lg_w_lg_w_q_range2333w2336w2337w2338w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_rad_ff2c_w_q_range2333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff3c	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff3c_w_lg_w_lg_w_q_range2365w2368w2369w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_rad_ff3c_w_lg_w_q_range2365w2366w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_rad_ff3c_w_lg_w_q_range2365w2368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff3c_w_lg_w_lg_w_lg_w_q_range2365w2368w2369w2370w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_rad_ff3c_w_q_range2365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff4c	:	STD_LOGIC_VECTOR(21 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff4c_w_lg_w_lg_w_q_range2397w2400w2401w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_rad_ff4c_w_lg_w_q_range2397w2398w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_rad_ff4c_w_lg_w_q_range2397w2400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff4c_w_lg_w_lg_w_lg_w_q_range2397w2400w2401w2402w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_rad_ff4c_w_q_range2397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff5c	:	STD_LOGIC_VECTOR(20 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff5c_w_lg_w_lg_w_q_range2429w2432w2433w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_rad_ff5c_w_lg_w_q_range2429w2430w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_rad_ff5c_w_lg_w_q_range2429w2432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff5c_w_lg_w_lg_w_lg_w_q_range2429w2432w2433w2434w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_rad_ff5c_w_q_range2429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff6c	:	STD_LOGIC_VECTOR(19 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff6c_w_lg_w_lg_w_q_range2461w2464w2465w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_rad_ff6c_w_lg_w_q_range2461w2462w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_rad_ff6c_w_lg_w_q_range2461w2464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff6c_w_lg_w_lg_w_lg_w_q_range2461w2464w2465w2466w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_rad_ff6c_w_q_range2461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff7c	:	STD_LOGIC_VECTOR(18 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff7c_w_lg_w_lg_w_q_range2493w2496w2497w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rad_ff7c_w_lg_w_q_range2493w2494w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rad_ff7c_w_lg_w_q_range2493w2496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff7c_w_lg_w_lg_w_lg_w_q_range2493w2496w2497w2498w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rad_ff7c_w_q_range2493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff8c	:	STD_LOGIC_VECTOR(17 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff8c_w_lg_w_lg_w_q_range2525w2528w2529w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_rad_ff8c_w_lg_w_q_range2525w2526w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_rad_ff8c_w_lg_w_q_range2525w2528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff8c_w_lg_w_lg_w_lg_w_q_range2525w2528w2529w2530w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_rad_ff8c_w_q_range2525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff9c	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff9c_w_lg_w_lg_w_q_range2557w2560w2561w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_rad_ff9c_w_lg_w_q_range2557w2558w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_rad_ff9c_w_lg_w_q_range2557w2560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff9c_w_lg_w_lg_w_lg_w_q_range2557w2560w2561w2562w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_rad_ff9c_w_q_range2557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub10_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub10_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub10_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub11_dataa	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_add_sub11_datab	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_add_sub11_result	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_add_sub12_dataa	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_add_sub12_datab	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_add_sub12_result	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_add_sub13_dataa	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub13_datab	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub13_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub14_dataa	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_add_sub14_datab	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_add_sub14_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_add_sub15_dataa	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_add_sub15_datab	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_add_sub15_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_add_sub16_dataa	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_add_sub16_datab	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_add_sub16_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_add_sub17_dataa	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_add_sub17_datab	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_add_sub17_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_add_sub18_dataa	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_add_sub18_datab	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_add_sub18_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_add_sub19_dataa	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_add_sub19_datab	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_add_sub19_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_add_sub20_dataa	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_add_sub20_datab	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_add_sub20_result	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_add_sub21_dataa	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_add_sub21_datab	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_add_sub21_result	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_add_sub22_dataa	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_add_sub22_datab	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_add_sub22_result	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_add_sub23_dataa	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_add_sub23_datab	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_add_sub23_result	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_add_sub24_dataa	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_add_sub24_datab	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_add_sub24_result	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_add_sub25_dataa	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_add_sub25_datab	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_add_sub25_result	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_add_sub26_dataa	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_add_sub26_datab	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_add_sub26_result	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_add_sub27_dataa	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_add_sub27_datab	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_add_sub27_result	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_add_sub28_dataa	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_add_sub28_datab	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_add_sub28_result	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_add_sub4_dataa	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_add_sub4_datab	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_add_sub4_result	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_add_sub5_dataa	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub5_datab	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub5_result	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub6_dataa	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_add_sub6_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_add_sub6_result	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_add_sub7_dataa	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_add_sub7_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_add_sub7_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_add_sub8_dataa	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_add_sub8_datab	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_add_sub8_result	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_add_sub9_dataa	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub9_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub9_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w10c_range914w915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w11c_range987w988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w12c_range1060w1061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w13c_range1133w1134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w14c_range1204w1205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w15c_range1275w1276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w16c_range1346w1347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w17c_range1417w1418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w18c_range1488w1489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w19c_range1559w1560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w1c_range257w258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w20c_range1630w1631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w21c_range1701w1702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w22c_range1772w1773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w23c_range1843w1844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w24c_range1914w1915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w2c_range330w331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w3c_range403w404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w4c_range476w477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w5c_range549w550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w6c_range622w623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w7c_range695w696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w8c_range768w769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w9c_range841w842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w10c_range2556w2559w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w11c_range2588w2591w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w12c_range2619w2622w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w13c_range2651w2654w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w14c_range2690w2693w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w15c_range2729w2732w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w16c_range2768w2771w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w17c_range2807w2810w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w18c_range2846w2849w	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w19c_range2885w2888w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w20c_range2924w2927w	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w21c_range2963w2966w	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w22c_range3002w3005w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w23c_range3041w3044w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w24c_range3083w3085w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w2c_range2300w2303w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w3c_range2332w2335w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w4c_range2364w2367w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w5c_range2396w2399w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w6c_range2428w2431w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w7c_range2460w2463w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w8c_range2492w2495w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w9c_range2524w2527w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  addnode_w0c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w10c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w11c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w12c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w13c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w14c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w15c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w16c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w17c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w18c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w19c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w1c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w20c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w21c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w22c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w23c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w24c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w2c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w3c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w4c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w5c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w6c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w7c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w8c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  addnode_w9c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  qlevel_w0c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  qlevel_w10c :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  qlevel_w11c :	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  qlevel_w12c :	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  qlevel_w13c :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  qlevel_w14c :	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  qlevel_w15c :	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  qlevel_w16c :	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  qlevel_w17c :	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  qlevel_w18c :	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  qlevel_w19c :	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  qlevel_w1c :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  qlevel_w20c :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  qlevel_w21c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  qlevel_w22c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  qlevel_w23c :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  qlevel_w24c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  qlevel_w2c :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  qlevel_w3c :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  qlevel_w4c :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  qlevel_w5c :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  qlevel_w6c :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  qlevel_w7c :	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  qlevel_w8c :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  qlevel_w9c :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  slevel_w0c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w10c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w11c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w12c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w13c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w14c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w15c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w16c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w17c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w18c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w19c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w1c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w20c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w21c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w22c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w23c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w24c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w2c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w3c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w4c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w5c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w6c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w7c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w8c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  slevel_w9c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w0c_range233w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w10c_range243w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w10c_range914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w11c_range244w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w11c_range987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w12c_range245w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w12c_range1060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w13c_range246w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w13c_range1133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w14c_range247w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w14c_range1204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w15c_range248w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w15c_range1275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w16c_range249w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w16c_range1346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w17c_range250w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w17c_range1417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w18c_range1488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w18c_range251w	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w19c_range1559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w19c_range252w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w1c_range234w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w1c_range257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w20c_range1630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w20c_range253w	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w21c_range1701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w21c_range254w	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w22c_range1772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w22c_range255w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w23c_range1843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w23c_range256w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w24c_range1914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w2c_range330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w2c_range235w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w3c_range403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w3c_range236w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w4c_range476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w4c_range237w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w5c_range549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w5c_range238w	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w6c_range622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w6c_range239w	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w7c_range695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w7c_range240w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w8c_range768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w8c_range241w	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w9c_range242w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w9c_range841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w10c_range2556w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w11c_range2588w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w12c_range2619w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w13c_range2651w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w14c_range2690w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w15c_range2729w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w16c_range2768w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w17c_range2807w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w18c_range2846w	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w19c_range2885w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w20c_range2924w	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w21c_range2963w	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w22c_range3002w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w23c_range3041w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w24c_range3083w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w2c_range2300w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w3c_range2332w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w4c_range2364w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w5c_range2396w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w6c_range2428w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w7c_range2460w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w8c_range2492w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w9c_range2524w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_alt_sqrt_block2_w_lg_w_addnode_w10c_range914w915w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w10c_range914w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w11c_range987w988w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w11c_range987w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w12c_range1060w1061w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w12c_range1060w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w13c_range1133w1134w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w13c_range1133w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w14c_range1204w1205w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w14c_range1204w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w15c_range1275w1276w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w15c_range1275w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w16c_range1346w1347w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w16c_range1346w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w17c_range1417w1418w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w17c_range1417w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w18c_range1488w1489w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w18c_range1488w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w19c_range1559w1560w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w19c_range1559w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w1c_range257w258w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w1c_range257w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w20c_range1630w1631w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w20c_range1630w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w21c_range1701w1702w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w21c_range1701w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w22c_range1772w1773w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w22c_range1772w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w23c_range1843w1844w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w23c_range1843w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w24c_range1914w1915w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w24c_range1914w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w2c_range330w331w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w2c_range330w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w3c_range403w404w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w3c_range403w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w4c_range476w477w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w4c_range476w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w5c_range549w550w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w5c_range549w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w6c_range622w623w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w6c_range622w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w7c_range695w696w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w7c_range695w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w8c_range768w769w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w8c_range768w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w9c_range841w842w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w9c_range841w(0);
	loop0 : FOR i IN 0 TO 10 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w10c_range2556w2559w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w10c_range2556w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 11 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w11c_range2588w2591w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w11c_range2588w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 12 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w12c_range2619w2622w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w12c_range2619w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 12 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w13c_range2651w2654w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w13c_range2651w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 13 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w14c_range2690w2693w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w14c_range2690w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 14 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w15c_range2729w2732w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w15c_range2729w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 15 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w16c_range2768w2771w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w16c_range2768w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 16 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w17c_range2807w2810w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w17c_range2807w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 17 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w18c_range2846w2849w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w18c_range2846w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 18 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w19c_range2885w2888w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w19c_range2885w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 19 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w20c_range2924w2927w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w20c_range2924w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 20 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w21c_range2963w2966w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w21c_range2963w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 21 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w22c_range3002w3005w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w22c_range3002w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 22 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w23c_range3041w3044w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w23c_range3041w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 21 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w24c_range3083w3085w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w24c_range3083w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 2 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w2c_range2300w2303w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w2c_range2300w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 3 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w3c_range2332w2335w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w3c_range2332w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 4 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w4c_range2364w2367w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w4c_range2364w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 5 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w5c_range2396w2399w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w5c_range2396w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 6 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w6c_range2428w2431w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w6c_range2428w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 7 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w7c_range2460w2463w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w7c_range2460w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 8 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w8c_range2492w2495w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w8c_range2492w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 9 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w9c_range2524w2527w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w9c_range2524w(i);
	END GENERATE loop22;
	addnode_w0c <= ( wire_add_sub4_result(2 DOWNTO 0) & slevel_w0c(23 DOWNTO 0));
	addnode_w10c <= ( wire_add_sub14_result(12 DOWNTO 0) & slevel_w10c(13 DOWNTO 0));
	addnode_w11c <= ( wire_add_sub15_result(13 DOWNTO 0) & slevel_w11c(12 DOWNTO 0));
	addnode_w12c <= ( wire_add_sub16_result(13 DOWNTO 0) & qlevel_w12c(0) & slevel_w12c(11 DOWNTO 0));
	addnode_w13c <= ( wire_add_sub17_result(12 DOWNTO 0) & "1" & qlevel_w13c(1 DOWNTO 0) & slevel_w13c(10 DOWNTO 0));
	addnode_w14c <= ( wire_add_sub18_result(13 DOWNTO 0) & "1" & qlevel_w14c(1 DOWNTO 0) & slevel_w14c(9 DOWNTO 0));
	addnode_w15c <= ( wire_add_sub19_result(14 DOWNTO 0) & "1" & qlevel_w15c(1 DOWNTO 0) & slevel_w15c(8 DOWNTO 0));
	addnode_w16c <= ( wire_add_sub20_result(15 DOWNTO 0) & "1" & qlevel_w16c(1 DOWNTO 0) & slevel_w16c(7 DOWNTO 0));
	addnode_w17c <= ( wire_add_sub21_result(16 DOWNTO 0) & "1" & qlevel_w17c(1 DOWNTO 0) & slevel_w17c(6 DOWNTO 0));
	addnode_w18c <= ( wire_add_sub22_result(17 DOWNTO 0) & "1" & qlevel_w18c(1 DOWNTO 0) & slevel_w18c(5 DOWNTO 0));
	addnode_w19c <= ( wire_add_sub23_result(18 DOWNTO 0) & "1" & qlevel_w19c(1 DOWNTO 0) & slevel_w19c(4 DOWNTO 0));
	addnode_w1c <= ( wire_add_sub5_result(3 DOWNTO 0) & slevel_w1c(22 DOWNTO 0));
	addnode_w20c <= ( wire_add_sub24_result(19 DOWNTO 0) & "1" & qlevel_w20c(1 DOWNTO 0) & slevel_w20c(3 DOWNTO 0));
	addnode_w21c <= ( wire_add_sub25_result(20 DOWNTO 0) & "1" & qlevel_w21c(1 DOWNTO 0) & slevel_w21c(2 DOWNTO 0));
	addnode_w22c <= ( wire_add_sub26_result(21 DOWNTO 0) & "1" & qlevel_w22c(1 DOWNTO 0) & slevel_w22c(1 DOWNTO 0));
	addnode_w23c <= ( wire_add_sub27_result(22 DOWNTO 0) & "1" & qlevel_w23c(1 DOWNTO 0) & slevel_w23c(0));
	addnode_w24c <= ( wire_add_sub28_result(23 DOWNTO 0) & "1" & qlevel_w24c(1 DOWNTO 0));
	addnode_w2c <= ( wire_add_sub6_result(4 DOWNTO 0) & slevel_w2c(21 DOWNTO 0));
	addnode_w3c <= ( wire_add_sub7_result(5 DOWNTO 0) & slevel_w3c(20 DOWNTO 0));
	addnode_w4c <= ( wire_add_sub8_result(6 DOWNTO 0) & slevel_w4c(19 DOWNTO 0));
	addnode_w5c <= ( wire_add_sub9_result(7 DOWNTO 0) & slevel_w5c(18 DOWNTO 0));
	addnode_w6c <= ( wire_add_sub10_result(8 DOWNTO 0) & slevel_w6c(17 DOWNTO 0));
	addnode_w7c <= ( wire_add_sub11_result(9 DOWNTO 0) & slevel_w7c(16 DOWNTO 0));
	addnode_w8c <= ( wire_add_sub12_result(10 DOWNTO 0) & slevel_w8c(15 DOWNTO 0));
	addnode_w9c <= ( wire_add_sub13_result(11 DOWNTO 0) & slevel_w9c(14 DOWNTO 0));
	qlevel_w0c <= ( "1" & "1" & "1");
	qlevel_w10c <= ( "0" & "1" & q_ff23c(8) & q_ff22c(7) & q_ff21c(6) & q_ff20c(5) & q_ff19c(4) & q_ff18c(3) & q_ff17c(2) & q_ff16c(1) & q_ff15c(0) & "1" & "1");
	qlevel_w11c <= ( "0" & "1" & q_ff23c(9) & q_ff22c(8) & q_ff21c(7) & q_ff20c(6) & q_ff19c(5) & q_ff18c(4) & q_ff17c(3) & q_ff16c(2) & q_ff15c(1) & q_ff14c(0) & "1" & "1");
	qlevel_w12c <= ( "0" & "1" & q_ff23c(10) & q_ff22c(9) & q_ff21c(8) & q_ff20c(7) & q_ff19c(6) & q_ff18c(5) & q_ff17c(4) & q_ff16c(3) & q_ff15c(2) & q_ff14c(1) & q_ff13c(0) & "1" & "1");
	qlevel_w13c <= ( "0" & "1" & q_ff23c(11) & q_ff22c(10) & q_ff21c(9) & q_ff20c(8) & q_ff19c(7) & q_ff18c(6) & q_ff17c(5) & q_ff16c(4) & q_ff15c(3) & q_ff14c(2) & q_ff13c(1) & q_ff12c(0) & "1" & "1");
	qlevel_w14c <= ( "0" & "1" & q_ff23c(12) & q_ff22c(11) & q_ff21c(10) & q_ff20c(9) & q_ff19c(8) & q_ff18c(7) & q_ff17c(6) & q_ff16c(5) & q_ff15c(4) & q_ff14c(3) & q_ff13c(2) & q_ff12c(1) & q_ff11c(0) & "1" & "1");
	qlevel_w15c <= ( "0" & "1" & q_ff23c(13) & q_ff22c(12) & q_ff21c(11) & q_ff20c(10) & q_ff19c(9) & q_ff18c(8) & q_ff17c(7) & q_ff16c(6) & q_ff15c(5) & q_ff14c(4) & q_ff13c(3) & q_ff12c(2) & q_ff11c(1) & q_ff10c(0) & "1" & "1");
	qlevel_w16c <= ( "0" & "1" & q_ff23c(14) & q_ff22c(13) & q_ff21c(12) & q_ff20c(11) & q_ff19c(10) & q_ff18c(9) & q_ff17c(8) & q_ff16c(7) & q_ff15c(6) & q_ff14c(5) & q_ff13c(4) & q_ff12c(3) & q_ff11c(2) & q_ff10c(1) & q_ff9c(0) & "1" & "1");
	qlevel_w17c <= ( "0" & "1" & q_ff23c(15) & q_ff22c(14) & q_ff21c(13) & q_ff20c(12) & q_ff19c(11) & q_ff18c(10) & q_ff17c(9) & q_ff16c(8) & q_ff15c(7) & q_ff14c(6) & q_ff13c(5) & q_ff12c(4) & q_ff11c(3) & q_ff10c(2) & q_ff9c(1) & q_ff8c(0) & "1" & "1");
	qlevel_w18c <= ( "0" & "1" & q_ff23c(16) & q_ff22c(15) & q_ff21c(14) & q_ff20c(13) & q_ff19c(12) & q_ff18c(11) & q_ff17c(10) & q_ff16c(9) & q_ff15c(8) & q_ff14c(7) & q_ff13c(6) & q_ff12c(5) & q_ff11c(4) & q_ff10c(3) & q_ff9c(2) & q_ff8c(1) & q_ff7c(0) & "1" & "1");
	qlevel_w19c <= ( "0" & "1" & q_ff23c(17) & q_ff22c(16) & q_ff21c(15) & q_ff20c(14) & q_ff19c(13) & q_ff18c(12) & q_ff17c(11) & q_ff16c(10) & q_ff15c(9) & q_ff14c(8) & q_ff13c(7) & q_ff12c(6) & q_ff11c(5) & q_ff10c(4) & q_ff9c(3) & q_ff8c(2) & q_ff7c(1) & q_ff6c(0) & "1" & "1");
	qlevel_w1c <= ( "1" & "0" & "1" & "1");
	qlevel_w20c <= ( "0" & "1" & q_ff23c(18) & q_ff22c(17) & q_ff21c(16) & q_ff20c(15) & q_ff19c(14) & q_ff18c(13) & q_ff17c(12) & q_ff16c(11) & q_ff15c(10) & q_ff14c(9) & q_ff13c(8) & q_ff12c(7) & q_ff11c(6) & q_ff10c(5) & q_ff9c(4) & q_ff8c(3) & q_ff7c(2) & q_ff6c(1) & q_ff5c(0) & "1" & "1");
	qlevel_w21c <= ( "0" & "1" & q_ff23c(19) & q_ff22c(18) & q_ff21c(17) & q_ff20c(16) & q_ff19c(15) & q_ff18c(14) & q_ff17c(13) & q_ff16c(12) & q_ff15c(11) & q_ff14c(10) & q_ff13c(9) & q_ff12c(8) & q_ff11c(7) & q_ff10c(6) & q_ff9c(5) & q_ff8c(4) & q_ff7c(3) & q_ff6c(2) & q_ff5c(1) & q_ff4c(0) & "1" & "1");
	qlevel_w22c <= ( "0" & "1" & q_ff23c(20) & q_ff22c(19) & q_ff21c(18) & q_ff20c(17) & q_ff19c(16) & q_ff18c(15) & q_ff17c(14) & q_ff16c(13) & q_ff15c(12) & q_ff14c(11) & q_ff13c(10) & q_ff12c(9) & q_ff11c(8) & q_ff10c(7) & q_ff9c(6) & q_ff8c(5) & q_ff7c(4) & q_ff6c(3) & q_ff5c(2) & q_ff4c(1) & q_ff3c(0) & "1" & "1");
	qlevel_w23c <= ( "0" & "1" & q_ff23c(21) & q_ff22c(20) & q_ff21c(19) & q_ff20c(18) & q_ff19c(17) & q_ff18c(16) & q_ff17c(15) & q_ff16c(14) & q_ff15c(13) & q_ff14c(12) & q_ff13c(11) & q_ff12c(10) & q_ff11c(9) & q_ff10c(8) & q_ff9c(7) & q_ff8c(6) & q_ff7c(5) & q_ff6c(4) & q_ff5c(3) & q_ff4c(2) & q_ff3c(1) & q_ff2c(0) & "1" & "1");
	qlevel_w24c <= ( wire_rad_ff23c_w_lg_w_q_range3069w3070w & rad_ff23c(22) & q_ff23c(22) & q_ff22c(21) & q_ff21c(20) & q_ff20c(19) & q_ff19c(18) & q_ff18c(17) & q_ff17c(16) & q_ff16c(15) & q_ff15c(14) & q_ff14c(13) & q_ff13c(12) & q_ff12c(11) & q_ff11c(10) & q_ff10c(9) & q_ff9c(8) & q_ff8c(7) & q_ff7c(6) & q_ff6c(5) & q_ff5c(4) & q_ff4c(3) & q_ff3c(2) & q_ff2c(1) & q_ff1c(0) & "1" & "1");
	qlevel_w2c <= ( "0" & "1" & q_ff23c(0) & "1" & "1");
	qlevel_w3c <= ( "0" & "1" & q_ff23c(1) & q_ff22c(0) & "1" & "1");
	qlevel_w4c <= ( "0" & "1" & q_ff23c(2) & q_ff22c(1) & q_ff21c(0) & "1" & "1");
	qlevel_w5c <= ( "0" & "1" & q_ff23c(3) & q_ff22c(2) & q_ff21c(1) & q_ff20c(0) & "1" & "1");
	qlevel_w6c <= ( "0" & "1" & q_ff23c(4) & q_ff22c(3) & q_ff21c(2) & q_ff20c(1) & q_ff19c(0) & "1" & "1");
	qlevel_w7c <= ( "0" & "1" & q_ff23c(5) & q_ff22c(4) & q_ff21c(3) & q_ff20c(2) & q_ff19c(1) & q_ff18c(0) & "1" & "1");
	qlevel_w8c <= ( "0" & "1" & q_ff23c(6) & q_ff22c(5) & q_ff21c(4) & q_ff20c(3) & q_ff19c(2) & q_ff18c(1) & q_ff17c(0) & "1" & "1");
	qlevel_w9c <= ( "0" & "1" & q_ff23c(7) & q_ff22c(6) & q_ff21c(5) & q_ff20c(4) & q_ff19c(3) & q_ff18c(2) & q_ff17c(1) & q_ff16c(0) & "1" & "1");
	root_result <= ( "1" & q_ff23c(23) & q_ff22c(22) & q_ff21c(21) & q_ff20c(20) & q_ff19c(19) & q_ff18c(18) & q_ff17c(17) & q_ff16c(16) & q_ff15c(15) & q_ff14c(14) & q_ff13c(13) & q_ff12c(12) & q_ff11c(11) & q_ff10c(10) & q_ff9c(9) & q_ff8c(8) & q_ff7c(7) & q_ff6c(6) & q_ff5c(5) & q_ff4c(4) & q_ff3c(3) & q_ff2c(2) & q_ff1c(1) & q_ff0c(0));
	slevel_w0c <= ( "0" & rad);
	slevel_w10c <= ( rad_ff9c(15 DOWNTO 0) & "00000000000");
	slevel_w11c <= ( rad_ff10c(14 DOWNTO 0) & "000000000000");
	slevel_w12c <= ( rad_ff11c(13 DOWNTO 0) & "0000000000000");
	slevel_w13c <= ( rad_ff12c(12 DOWNTO 0) & "1" & "0000000000000");
	slevel_w14c <= ( rad_ff13c(11 DOWNTO 0) & "1" & "1" & "1" & "000000000000");
	slevel_w15c <= ( rad_ff14c(12 DOWNTO 0) & "1" & "1" & "1" & "00000000000");
	slevel_w16c <= ( rad_ff15c(13 DOWNTO 0) & "1" & "1" & "1" & "0000000000");
	slevel_w17c <= ( rad_ff16c(14 DOWNTO 0) & "1" & "1" & "1" & "000000000");
	slevel_w18c <= ( rad_ff17c(15 DOWNTO 0) & "1" & "1" & "1" & "00000000");
	slevel_w19c <= ( rad_ff18c(16 DOWNTO 0) & "1" & "1" & "1" & "0000000");
	slevel_w1c <= ( rad_ff0c(24 DOWNTO 0) & "0" & "0");
	slevel_w20c <= ( rad_ff19c(17 DOWNTO 0) & "1" & "1" & "1" & "000000");
	slevel_w21c <= ( rad_ff20c(18 DOWNTO 0) & "1" & "1" & "1" & "00000");
	slevel_w22c <= ( rad_ff21c(19 DOWNTO 0) & "1" & "1" & "1" & "0000");
	slevel_w23c <= ( rad_ff22c(20 DOWNTO 0) & "1" & "1" & "1" & "000");
	slevel_w24c <= ( rad_ff23c(21 DOWNTO 0) & "1" & "1" & "1" & "00");
	slevel_w2c <= ( rad_ff1c(23 DOWNTO 0) & "000");
	slevel_w3c <= ( rad_ff2c(22 DOWNTO 0) & "0000");
	slevel_w4c <= ( rad_ff3c(21 DOWNTO 0) & "00000");
	slevel_w5c <= ( rad_ff4c(20 DOWNTO 0) & "000000");
	slevel_w6c <= ( rad_ff5c(19 DOWNTO 0) & "0000000");
	slevel_w7c <= ( rad_ff6c(18 DOWNTO 0) & "00000000");
	slevel_w8c <= ( rad_ff7c(17 DOWNTO 0) & "000000000");
	slevel_w9c <= ( rad_ff8c(16 DOWNTO 0) & "0000000000");
	wire_alt_sqrt_block2_w_addnode_w0c_range233w <= addnode_w0c(26 DOWNTO 1);
	wire_alt_sqrt_block2_w_addnode_w10c_range243w <= addnode_w10c(26 DOWNTO 11);
	wire_alt_sqrt_block2_w_addnode_w10c_range914w(0) <= addnode_w10c(26);
	wire_alt_sqrt_block2_w_addnode_w11c_range244w <= addnode_w11c(26 DOWNTO 12);
	wire_alt_sqrt_block2_w_addnode_w11c_range987w(0) <= addnode_w11c(26);
	wire_alt_sqrt_block2_w_addnode_w12c_range245w <= addnode_w12c(26 DOWNTO 13);
	wire_alt_sqrt_block2_w_addnode_w12c_range1060w(0) <= addnode_w12c(26);
	wire_alt_sqrt_block2_w_addnode_w13c_range246w <= addnode_w13c(26 DOWNTO 14);
	wire_alt_sqrt_block2_w_addnode_w13c_range1133w(0) <= addnode_w13c(26);
	wire_alt_sqrt_block2_w_addnode_w14c_range247w <= addnode_w14c(26 DOWNTO 13);
	wire_alt_sqrt_block2_w_addnode_w14c_range1204w(0) <= addnode_w14c(26);
	wire_alt_sqrt_block2_w_addnode_w15c_range248w <= addnode_w15c(26 DOWNTO 12);
	wire_alt_sqrt_block2_w_addnode_w15c_range1275w(0) <= addnode_w15c(26);
	wire_alt_sqrt_block2_w_addnode_w16c_range249w <= addnode_w16c(26 DOWNTO 11);
	wire_alt_sqrt_block2_w_addnode_w16c_range1346w(0) <= addnode_w16c(26);
	wire_alt_sqrt_block2_w_addnode_w17c_range250w <= addnode_w17c(26 DOWNTO 10);
	wire_alt_sqrt_block2_w_addnode_w17c_range1417w(0) <= addnode_w17c(26);
	wire_alt_sqrt_block2_w_addnode_w18c_range1488w(0) <= addnode_w18c(26);
	wire_alt_sqrt_block2_w_addnode_w18c_range251w <= addnode_w18c(26 DOWNTO 9);
	wire_alt_sqrt_block2_w_addnode_w19c_range1559w(0) <= addnode_w19c(26);
	wire_alt_sqrt_block2_w_addnode_w19c_range252w <= addnode_w19c(26 DOWNTO 8);
	wire_alt_sqrt_block2_w_addnode_w1c_range234w <= addnode_w1c(26 DOWNTO 2);
	wire_alt_sqrt_block2_w_addnode_w1c_range257w(0) <= addnode_w1c(26);
	wire_alt_sqrt_block2_w_addnode_w20c_range1630w(0) <= addnode_w20c(26);
	wire_alt_sqrt_block2_w_addnode_w20c_range253w <= addnode_w20c(26 DOWNTO 7);
	wire_alt_sqrt_block2_w_addnode_w21c_range1701w(0) <= addnode_w21c(26);
	wire_alt_sqrt_block2_w_addnode_w21c_range254w <= addnode_w21c(26 DOWNTO 6);
	wire_alt_sqrt_block2_w_addnode_w22c_range1772w(0) <= addnode_w22c(26);
	wire_alt_sqrt_block2_w_addnode_w22c_range255w <= addnode_w22c(26 DOWNTO 5);
	wire_alt_sqrt_block2_w_addnode_w23c_range1843w(0) <= addnode_w23c(26);
	wire_alt_sqrt_block2_w_addnode_w23c_range256w <= addnode_w23c(26 DOWNTO 4);
	wire_alt_sqrt_block2_w_addnode_w24c_range1914w(0) <= addnode_w24c(26);
	wire_alt_sqrt_block2_w_addnode_w2c_range330w(0) <= addnode_w2c(26);
	wire_alt_sqrt_block2_w_addnode_w2c_range235w <= addnode_w2c(26 DOWNTO 3);
	wire_alt_sqrt_block2_w_addnode_w3c_range403w(0) <= addnode_w3c(26);
	wire_alt_sqrt_block2_w_addnode_w3c_range236w <= addnode_w3c(26 DOWNTO 4);
	wire_alt_sqrt_block2_w_addnode_w4c_range476w(0) <= addnode_w4c(26);
	wire_alt_sqrt_block2_w_addnode_w4c_range237w <= addnode_w4c(26 DOWNTO 5);
	wire_alt_sqrt_block2_w_addnode_w5c_range549w(0) <= addnode_w5c(26);
	wire_alt_sqrt_block2_w_addnode_w5c_range238w <= addnode_w5c(26 DOWNTO 6);
	wire_alt_sqrt_block2_w_addnode_w6c_range622w(0) <= addnode_w6c(26);
	wire_alt_sqrt_block2_w_addnode_w6c_range239w <= addnode_w6c(26 DOWNTO 7);
	wire_alt_sqrt_block2_w_addnode_w7c_range695w(0) <= addnode_w7c(26);
	wire_alt_sqrt_block2_w_addnode_w7c_range240w <= addnode_w7c(26 DOWNTO 8);
	wire_alt_sqrt_block2_w_addnode_w8c_range768w(0) <= addnode_w8c(26);
	wire_alt_sqrt_block2_w_addnode_w8c_range241w <= addnode_w8c(26 DOWNTO 9);
	wire_alt_sqrt_block2_w_addnode_w9c_range242w <= addnode_w9c(26 DOWNTO 10);
	wire_alt_sqrt_block2_w_addnode_w9c_range841w(0) <= addnode_w9c(26);
	wire_alt_sqrt_block2_w_qlevel_w10c_range2556w <= qlevel_w10c(12 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w11c_range2588w <= qlevel_w11c(13 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w12c_range2619w <= qlevel_w12c(14 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w13c_range2651w <= qlevel_w13c(15 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w14c_range2690w <= qlevel_w14c(16 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w15c_range2729w <= qlevel_w15c(17 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w16c_range2768w <= qlevel_w16c(18 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w17c_range2807w <= qlevel_w17c(19 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w18c_range2846w <= qlevel_w18c(20 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w19c_range2885w <= qlevel_w19c(21 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w20c_range2924w <= qlevel_w20c(22 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w21c_range2963w <= qlevel_w21c(23 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w22c_range3002w <= qlevel_w22c(24 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w23c_range3041w <= qlevel_w23c(25 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w24c_range3083w <= qlevel_w24c(24 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w2c_range2300w <= qlevel_w2c(4 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w3c_range2332w <= qlevel_w3c(5 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w4c_range2364w <= qlevel_w4c(6 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w5c_range2396w <= qlevel_w5c(7 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w6c_range2428w <= qlevel_w6c(8 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w7c_range2460w <= qlevel_w7c(9 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w8c_range2492w <= qlevel_w8c(10 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w9c_range2524w <= qlevel_w9c(11 DOWNTO 2);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff0c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff0c <= ( q_ff0c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w24c_range1914w1915w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff10c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff10c <= ( q_ff10c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w14c_range1204w1205w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff11c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff11c <= ( q_ff11c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w13c_range1133w1134w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff12c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff12c <= ( q_ff12c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w12c_range1060w1061w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff13c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff13c <= ( q_ff13c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w11c_range987w988w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff14c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff14c <= ( q_ff14c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w10c_range914w915w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff15c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff15c <= ( q_ff15c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w9c_range841w842w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff16c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff16c <= ( q_ff16c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w8c_range768w769w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff17c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff17c <= ( q_ff17c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w7c_range695w696w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff18c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff18c <= ( q_ff18c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w6c_range622w623w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff19c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff19c <= ( q_ff19c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w5c_range549w550w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff1c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff1c <= ( q_ff1c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w23c_range1843w1844w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff20c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff20c <= ( q_ff20c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w4c_range476w477w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff21c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff21c <= ( q_ff21c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w3c_range403w404w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff22c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff22c <= ( q_ff22c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w2c_range330w331w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff23c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff23c <= ( q_ff23c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w1c_range257w258w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff2c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff2c <= ( q_ff2c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w22c_range1772w1773w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff3c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff3c <= ( q_ff3c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w21c_range1701w1702w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff4c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff4c <= ( q_ff4c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w20c_range1630w1631w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff5c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff5c <= ( q_ff5c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w19c_range1559w1560w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff6c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff6c <= ( q_ff6c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w18c_range1488w1489w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff7c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff7c <= ( q_ff7c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w17c_range1417w1418w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff8c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff8c <= ( q_ff8c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w16c_range1346w1347w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff9c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff9c <= ( q_ff9c(22 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w15c_range1275w1276w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff0c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff0c <= wire_alt_sqrt_block2_w_addnode_w0c_range233w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff10c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff10c <= wire_alt_sqrt_block2_w_addnode_w10c_range243w;
			END IF;
		END IF;
	END PROCESS;
	loop23 : FOR i IN 0 TO 11 GENERATE 
		wire_rad_ff10c_w_lg_w_lg_w_q_range2589w2592w2593w(i) <= wire_rad_ff10c_w_lg_w_q_range2589w2592w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w11c_range2588w2591w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 11 GENERATE 
		wire_rad_ff10c_w_lg_w_q_range2589w2590w(i) <= wire_rad_ff10c_w_q_range2589w(0) AND wire_alt_sqrt_block2_w_qlevel_w11c_range2588w(i);
	END GENERATE loop24;
	wire_rad_ff10c_w_lg_w_q_range2589w2592w(0) <= NOT wire_rad_ff10c_w_q_range2589w(0);
	loop25 : FOR i IN 0 TO 11 GENERATE 
		wire_rad_ff10c_w_lg_w_lg_w_lg_w_q_range2589w2592w2593w2594w(i) <= wire_rad_ff10c_w_lg_w_lg_w_q_range2589w2592w2593w(i) OR wire_rad_ff10c_w_lg_w_q_range2589w2590w(i);
	END GENERATE loop25;
	wire_rad_ff10c_w_q_range2589w(0) <= rad_ff10c(15);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff11c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff11c <= wire_alt_sqrt_block2_w_addnode_w11c_range244w;
			END IF;
		END IF;
	END PROCESS;
	loop26 : FOR i IN 0 TO 12 GENERATE 
		wire_rad_ff11c_w_lg_w_lg_w_q_range2620w2623w2624w(i) <= wire_rad_ff11c_w_lg_w_q_range2620w2623w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w12c_range2619w2622w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 12 GENERATE 
		wire_rad_ff11c_w_lg_w_q_range2620w2621w(i) <= wire_rad_ff11c_w_q_range2620w(0) AND wire_alt_sqrt_block2_w_qlevel_w12c_range2619w(i);
	END GENERATE loop27;
	wire_rad_ff11c_w_lg_w_q_range2620w2623w(0) <= NOT wire_rad_ff11c_w_q_range2620w(0);
	loop28 : FOR i IN 0 TO 12 GENERATE 
		wire_rad_ff11c_w_lg_w_lg_w_lg_w_q_range2620w2623w2624w2625w(i) <= wire_rad_ff11c_w_lg_w_lg_w_q_range2620w2623w2624w(i) OR wire_rad_ff11c_w_lg_w_q_range2620w2621w(i);
	END GENERATE loop28;
	wire_rad_ff11c_w_q_range2620w(0) <= rad_ff11c(14);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff12c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff12c <= wire_alt_sqrt_block2_w_addnode_w12c_range245w;
			END IF;
		END IF;
	END PROCESS;
	loop29 : FOR i IN 0 TO 12 GENERATE 
		wire_rad_ff12c_w_lg_w_lg_w_q_range2652w2655w2656w(i) <= wire_rad_ff12c_w_lg_w_q_range2652w2655w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w13c_range2651w2654w(i);
	END GENERATE loop29;
	loop30 : FOR i IN 0 TO 12 GENERATE 
		wire_rad_ff12c_w_lg_w_q_range2652w2653w(i) <= wire_rad_ff12c_w_q_range2652w(0) AND wire_alt_sqrt_block2_w_qlevel_w13c_range2651w(i);
	END GENERATE loop30;
	wire_rad_ff12c_w_lg_w_q_range2652w2655w(0) <= NOT wire_rad_ff12c_w_q_range2652w(0);
	loop31 : FOR i IN 0 TO 12 GENERATE 
		wire_rad_ff12c_w_lg_w_lg_w_lg_w_q_range2652w2655w2656w2657w(i) <= wire_rad_ff12c_w_lg_w_lg_w_q_range2652w2655w2656w(i) OR wire_rad_ff12c_w_lg_w_q_range2652w2653w(i);
	END GENERATE loop31;
	wire_rad_ff12c_w_q_range2652w(0) <= rad_ff12c(13);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff13c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff13c <= wire_alt_sqrt_block2_w_addnode_w13c_range246w;
			END IF;
		END IF;
	END PROCESS;
	loop32 : FOR i IN 0 TO 13 GENERATE 
		wire_rad_ff13c_w_lg_w_lg_w_q_range2691w2694w2695w(i) <= wire_rad_ff13c_w_lg_w_q_range2691w2694w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w14c_range2690w2693w(i);
	END GENERATE loop32;
	loop33 : FOR i IN 0 TO 13 GENERATE 
		wire_rad_ff13c_w_lg_w_q_range2691w2692w(i) <= wire_rad_ff13c_w_q_range2691w(0) AND wire_alt_sqrt_block2_w_qlevel_w14c_range2690w(i);
	END GENERATE loop33;
	wire_rad_ff13c_w_lg_w_q_range2691w2694w(0) <= NOT wire_rad_ff13c_w_q_range2691w(0);
	loop34 : FOR i IN 0 TO 13 GENERATE 
		wire_rad_ff13c_w_lg_w_lg_w_lg_w_q_range2691w2694w2695w2696w(i) <= wire_rad_ff13c_w_lg_w_lg_w_q_range2691w2694w2695w(i) OR wire_rad_ff13c_w_lg_w_q_range2691w2692w(i);
	END GENERATE loop34;
	wire_rad_ff13c_w_q_range2691w(0) <= rad_ff13c(12);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff14c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff14c <= wire_alt_sqrt_block2_w_addnode_w14c_range247w;
			END IF;
		END IF;
	END PROCESS;
	loop35 : FOR i IN 0 TO 14 GENERATE 
		wire_rad_ff14c_w_lg_w_lg_w_q_range2730w2733w2734w(i) <= wire_rad_ff14c_w_lg_w_q_range2730w2733w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w15c_range2729w2732w(i);
	END GENERATE loop35;
	loop36 : FOR i IN 0 TO 14 GENERATE 
		wire_rad_ff14c_w_lg_w_q_range2730w2731w(i) <= wire_rad_ff14c_w_q_range2730w(0) AND wire_alt_sqrt_block2_w_qlevel_w15c_range2729w(i);
	END GENERATE loop36;
	wire_rad_ff14c_w_lg_w_q_range2730w2733w(0) <= NOT wire_rad_ff14c_w_q_range2730w(0);
	loop37 : FOR i IN 0 TO 14 GENERATE 
		wire_rad_ff14c_w_lg_w_lg_w_lg_w_q_range2730w2733w2734w2735w(i) <= wire_rad_ff14c_w_lg_w_lg_w_q_range2730w2733w2734w(i) OR wire_rad_ff14c_w_lg_w_q_range2730w2731w(i);
	END GENERATE loop37;
	wire_rad_ff14c_w_q_range2730w(0) <= rad_ff14c(13);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff15c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff15c <= wire_alt_sqrt_block2_w_addnode_w15c_range248w;
			END IF;
		END IF;
	END PROCESS;
	loop38 : FOR i IN 0 TO 15 GENERATE 
		wire_rad_ff15c_w_lg_w_lg_w_q_range2769w2772w2773w(i) <= wire_rad_ff15c_w_lg_w_q_range2769w2772w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w16c_range2768w2771w(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 15 GENERATE 
		wire_rad_ff15c_w_lg_w_q_range2769w2770w(i) <= wire_rad_ff15c_w_q_range2769w(0) AND wire_alt_sqrt_block2_w_qlevel_w16c_range2768w(i);
	END GENERATE loop39;
	wire_rad_ff15c_w_lg_w_q_range2769w2772w(0) <= NOT wire_rad_ff15c_w_q_range2769w(0);
	loop40 : FOR i IN 0 TO 15 GENERATE 
		wire_rad_ff15c_w_lg_w_lg_w_lg_w_q_range2769w2772w2773w2774w(i) <= wire_rad_ff15c_w_lg_w_lg_w_q_range2769w2772w2773w(i) OR wire_rad_ff15c_w_lg_w_q_range2769w2770w(i);
	END GENERATE loop40;
	wire_rad_ff15c_w_q_range2769w(0) <= rad_ff15c(14);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff16c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff16c <= wire_alt_sqrt_block2_w_addnode_w16c_range249w;
			END IF;
		END IF;
	END PROCESS;
	loop41 : FOR i IN 0 TO 16 GENERATE 
		wire_rad_ff16c_w_lg_w_lg_w_q_range2808w2811w2812w(i) <= wire_rad_ff16c_w_lg_w_q_range2808w2811w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w17c_range2807w2810w(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 16 GENERATE 
		wire_rad_ff16c_w_lg_w_q_range2808w2809w(i) <= wire_rad_ff16c_w_q_range2808w(0) AND wire_alt_sqrt_block2_w_qlevel_w17c_range2807w(i);
	END GENERATE loop42;
	wire_rad_ff16c_w_lg_w_q_range2808w2811w(0) <= NOT wire_rad_ff16c_w_q_range2808w(0);
	loop43 : FOR i IN 0 TO 16 GENERATE 
		wire_rad_ff16c_w_lg_w_lg_w_lg_w_q_range2808w2811w2812w2813w(i) <= wire_rad_ff16c_w_lg_w_lg_w_q_range2808w2811w2812w(i) OR wire_rad_ff16c_w_lg_w_q_range2808w2809w(i);
	END GENERATE loop43;
	wire_rad_ff16c_w_q_range2808w(0) <= rad_ff16c(15);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff17c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff17c <= wire_alt_sqrt_block2_w_addnode_w17c_range250w;
			END IF;
		END IF;
	END PROCESS;
	loop44 : FOR i IN 0 TO 17 GENERATE 
		wire_rad_ff17c_w_lg_w_lg_w_q_range2847w2850w2851w(i) <= wire_rad_ff17c_w_lg_w_q_range2847w2850w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w18c_range2846w2849w(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 17 GENERATE 
		wire_rad_ff17c_w_lg_w_q_range2847w2848w(i) <= wire_rad_ff17c_w_q_range2847w(0) AND wire_alt_sqrt_block2_w_qlevel_w18c_range2846w(i);
	END GENERATE loop45;
	wire_rad_ff17c_w_lg_w_q_range2847w2850w(0) <= NOT wire_rad_ff17c_w_q_range2847w(0);
	loop46 : FOR i IN 0 TO 17 GENERATE 
		wire_rad_ff17c_w_lg_w_lg_w_lg_w_q_range2847w2850w2851w2852w(i) <= wire_rad_ff17c_w_lg_w_lg_w_q_range2847w2850w2851w(i) OR wire_rad_ff17c_w_lg_w_q_range2847w2848w(i);
	END GENERATE loop46;
	wire_rad_ff17c_w_q_range2847w(0) <= rad_ff17c(16);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff18c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff18c <= wire_alt_sqrt_block2_w_addnode_w18c_range251w;
			END IF;
		END IF;
	END PROCESS;
	loop47 : FOR i IN 0 TO 18 GENERATE 
		wire_rad_ff18c_w_lg_w_lg_w_q_range2886w2889w2890w(i) <= wire_rad_ff18c_w_lg_w_q_range2886w2889w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w19c_range2885w2888w(i);
	END GENERATE loop47;
	loop48 : FOR i IN 0 TO 18 GENERATE 
		wire_rad_ff18c_w_lg_w_q_range2886w2887w(i) <= wire_rad_ff18c_w_q_range2886w(0) AND wire_alt_sqrt_block2_w_qlevel_w19c_range2885w(i);
	END GENERATE loop48;
	wire_rad_ff18c_w_lg_w_q_range2886w2889w(0) <= NOT wire_rad_ff18c_w_q_range2886w(0);
	loop49 : FOR i IN 0 TO 18 GENERATE 
		wire_rad_ff18c_w_lg_w_lg_w_lg_w_q_range2886w2889w2890w2891w(i) <= wire_rad_ff18c_w_lg_w_lg_w_q_range2886w2889w2890w(i) OR wire_rad_ff18c_w_lg_w_q_range2886w2887w(i);
	END GENERATE loop49;
	wire_rad_ff18c_w_q_range2886w(0) <= rad_ff18c(17);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff19c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff19c <= wire_alt_sqrt_block2_w_addnode_w19c_range252w;
			END IF;
		END IF;
	END PROCESS;
	loop50 : FOR i IN 0 TO 19 GENERATE 
		wire_rad_ff19c_w_lg_w_lg_w_q_range2925w2928w2929w(i) <= wire_rad_ff19c_w_lg_w_q_range2925w2928w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w20c_range2924w2927w(i);
	END GENERATE loop50;
	loop51 : FOR i IN 0 TO 19 GENERATE 
		wire_rad_ff19c_w_lg_w_q_range2925w2926w(i) <= wire_rad_ff19c_w_q_range2925w(0) AND wire_alt_sqrt_block2_w_qlevel_w20c_range2924w(i);
	END GENERATE loop51;
	wire_rad_ff19c_w_lg_w_q_range2925w2928w(0) <= NOT wire_rad_ff19c_w_q_range2925w(0);
	loop52 : FOR i IN 0 TO 19 GENERATE 
		wire_rad_ff19c_w_lg_w_lg_w_lg_w_q_range2925w2928w2929w2930w(i) <= wire_rad_ff19c_w_lg_w_lg_w_q_range2925w2928w2929w(i) OR wire_rad_ff19c_w_lg_w_q_range2925w2926w(i);
	END GENERATE loop52;
	wire_rad_ff19c_w_q_range2925w(0) <= rad_ff19c(18);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff1c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff1c <= wire_alt_sqrt_block2_w_addnode_w1c_range234w;
			END IF;
		END IF;
	END PROCESS;
	loop53 : FOR i IN 0 TO 2 GENERATE 
		wire_rad_ff1c_w_lg_w_lg_w_q_range2301w2304w2305w(i) <= wire_rad_ff1c_w_lg_w_q_range2301w2304w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w2c_range2300w2303w(i);
	END GENERATE loop53;
	loop54 : FOR i IN 0 TO 2 GENERATE 
		wire_rad_ff1c_w_lg_w_q_range2301w2302w(i) <= wire_rad_ff1c_w_q_range2301w(0) AND wire_alt_sqrt_block2_w_qlevel_w2c_range2300w(i);
	END GENERATE loop54;
	wire_rad_ff1c_w_lg_w_q_range2301w2304w(0) <= NOT wire_rad_ff1c_w_q_range2301w(0);
	loop55 : FOR i IN 0 TO 2 GENERATE 
		wire_rad_ff1c_w_lg_w_lg_w_lg_w_q_range2301w2304w2305w2306w(i) <= wire_rad_ff1c_w_lg_w_lg_w_q_range2301w2304w2305w(i) OR wire_rad_ff1c_w_lg_w_q_range2301w2302w(i);
	END GENERATE loop55;
	wire_rad_ff1c_w_q_range2301w(0) <= rad_ff1c(24);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff20c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff20c <= wire_alt_sqrt_block2_w_addnode_w20c_range253w;
			END IF;
		END IF;
	END PROCESS;
	loop56 : FOR i IN 0 TO 20 GENERATE 
		wire_rad_ff20c_w_lg_w_lg_w_q_range2964w2967w2968w(i) <= wire_rad_ff20c_w_lg_w_q_range2964w2967w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w21c_range2963w2966w(i);
	END GENERATE loop56;
	loop57 : FOR i IN 0 TO 20 GENERATE 
		wire_rad_ff20c_w_lg_w_q_range2964w2965w(i) <= wire_rad_ff20c_w_q_range2964w(0) AND wire_alt_sqrt_block2_w_qlevel_w21c_range2963w(i);
	END GENERATE loop57;
	wire_rad_ff20c_w_lg_w_q_range2964w2967w(0) <= NOT wire_rad_ff20c_w_q_range2964w(0);
	loop58 : FOR i IN 0 TO 20 GENERATE 
		wire_rad_ff20c_w_lg_w_lg_w_lg_w_q_range2964w2967w2968w2969w(i) <= wire_rad_ff20c_w_lg_w_lg_w_q_range2964w2967w2968w(i) OR wire_rad_ff20c_w_lg_w_q_range2964w2965w(i);
	END GENERATE loop58;
	wire_rad_ff20c_w_q_range2964w(0) <= rad_ff20c(19);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff21c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff21c <= wire_alt_sqrt_block2_w_addnode_w21c_range254w;
			END IF;
		END IF;
	END PROCESS;
	loop59 : FOR i IN 0 TO 21 GENERATE 
		wire_rad_ff21c_w_lg_w_lg_w_q_range3003w3006w3007w(i) <= wire_rad_ff21c_w_lg_w_q_range3003w3006w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w22c_range3002w3005w(i);
	END GENERATE loop59;
	loop60 : FOR i IN 0 TO 21 GENERATE 
		wire_rad_ff21c_w_lg_w_q_range3003w3004w(i) <= wire_rad_ff21c_w_q_range3003w(0) AND wire_alt_sqrt_block2_w_qlevel_w22c_range3002w(i);
	END GENERATE loop60;
	wire_rad_ff21c_w_lg_w_q_range3003w3006w(0) <= NOT wire_rad_ff21c_w_q_range3003w(0);
	loop61 : FOR i IN 0 TO 21 GENERATE 
		wire_rad_ff21c_w_lg_w_lg_w_lg_w_q_range3003w3006w3007w3008w(i) <= wire_rad_ff21c_w_lg_w_lg_w_q_range3003w3006w3007w(i) OR wire_rad_ff21c_w_lg_w_q_range3003w3004w(i);
	END GENERATE loop61;
	wire_rad_ff21c_w_q_range3003w(0) <= rad_ff21c(20);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff22c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff22c <= wire_alt_sqrt_block2_w_addnode_w22c_range255w;
			END IF;
		END IF;
	END PROCESS;
	loop62 : FOR i IN 0 TO 22 GENERATE 
		wire_rad_ff22c_w_lg_w_lg_w_q_range3042w3045w3046w(i) <= wire_rad_ff22c_w_lg_w_q_range3042w3045w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w23c_range3041w3044w(i);
	END GENERATE loop62;
	loop63 : FOR i IN 0 TO 22 GENERATE 
		wire_rad_ff22c_w_lg_w_q_range3042w3043w(i) <= wire_rad_ff22c_w_q_range3042w(0) AND wire_alt_sqrt_block2_w_qlevel_w23c_range3041w(i);
	END GENERATE loop63;
	wire_rad_ff22c_w_lg_w_q_range3042w3045w(0) <= NOT wire_rad_ff22c_w_q_range3042w(0);
	loop64 : FOR i IN 0 TO 22 GENERATE 
		wire_rad_ff22c_w_lg_w_lg_w_lg_w_q_range3042w3045w3046w3047w(i) <= wire_rad_ff22c_w_lg_w_lg_w_q_range3042w3045w3046w(i) OR wire_rad_ff22c_w_lg_w_q_range3042w3043w(i);
	END GENERATE loop64;
	wire_rad_ff22c_w_q_range3042w(0) <= rad_ff22c(21);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff23c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff23c <= wire_alt_sqrt_block2_w_addnode_w23c_range256w;
			END IF;
		END IF;
	END PROCESS;
	loop65 : FOR i IN 0 TO 21 GENERATE 
		wire_rad_ff23c_w_lg_w_lg_w_q_range3069w3070w3086w(i) <= wire_rad_ff23c_w_lg_w_q_range3069w3070w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w24c_range3083w3085w(i);
	END GENERATE loop65;
	loop66 : FOR i IN 0 TO 21 GENERATE 
		wire_rad_ff23c_w_lg_w_q_range3069w3084w(i) <= wire_rad_ff23c_w_q_range3069w(0) AND wire_alt_sqrt_block2_w_qlevel_w24c_range3083w(i);
	END GENERATE loop66;
	wire_rad_ff23c_w_lg_w_q_range3069w3070w(0) <= NOT wire_rad_ff23c_w_q_range3069w(0);
	loop67 : FOR i IN 0 TO 21 GENERATE 
		wire_rad_ff23c_w_lg_w_lg_w_lg_w_q_range3069w3070w3086w3087w(i) <= wire_rad_ff23c_w_lg_w_lg_w_q_range3069w3070w3086w(i) OR wire_rad_ff23c_w_lg_w_q_range3069w3084w(i);
	END GENERATE loop67;
	wire_rad_ff23c_w_q_range3069w(0) <= rad_ff23c(22);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff2c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff2c <= wire_alt_sqrt_block2_w_addnode_w2c_range235w;
			END IF;
		END IF;
	END PROCESS;
	loop68 : FOR i IN 0 TO 3 GENERATE 
		wire_rad_ff2c_w_lg_w_lg_w_q_range2333w2336w2337w(i) <= wire_rad_ff2c_w_lg_w_q_range2333w2336w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w3c_range2332w2335w(i);
	END GENERATE loop68;
	loop69 : FOR i IN 0 TO 3 GENERATE 
		wire_rad_ff2c_w_lg_w_q_range2333w2334w(i) <= wire_rad_ff2c_w_q_range2333w(0) AND wire_alt_sqrt_block2_w_qlevel_w3c_range2332w(i);
	END GENERATE loop69;
	wire_rad_ff2c_w_lg_w_q_range2333w2336w(0) <= NOT wire_rad_ff2c_w_q_range2333w(0);
	loop70 : FOR i IN 0 TO 3 GENERATE 
		wire_rad_ff2c_w_lg_w_lg_w_lg_w_q_range2333w2336w2337w2338w(i) <= wire_rad_ff2c_w_lg_w_lg_w_q_range2333w2336w2337w(i) OR wire_rad_ff2c_w_lg_w_q_range2333w2334w(i);
	END GENERATE loop70;
	wire_rad_ff2c_w_q_range2333w(0) <= rad_ff2c(23);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff3c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff3c <= wire_alt_sqrt_block2_w_addnode_w3c_range236w;
			END IF;
		END IF;
	END PROCESS;
	loop71 : FOR i IN 0 TO 4 GENERATE 
		wire_rad_ff3c_w_lg_w_lg_w_q_range2365w2368w2369w(i) <= wire_rad_ff3c_w_lg_w_q_range2365w2368w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w4c_range2364w2367w(i);
	END GENERATE loop71;
	loop72 : FOR i IN 0 TO 4 GENERATE 
		wire_rad_ff3c_w_lg_w_q_range2365w2366w(i) <= wire_rad_ff3c_w_q_range2365w(0) AND wire_alt_sqrt_block2_w_qlevel_w4c_range2364w(i);
	END GENERATE loop72;
	wire_rad_ff3c_w_lg_w_q_range2365w2368w(0) <= NOT wire_rad_ff3c_w_q_range2365w(0);
	loop73 : FOR i IN 0 TO 4 GENERATE 
		wire_rad_ff3c_w_lg_w_lg_w_lg_w_q_range2365w2368w2369w2370w(i) <= wire_rad_ff3c_w_lg_w_lg_w_q_range2365w2368w2369w(i) OR wire_rad_ff3c_w_lg_w_q_range2365w2366w(i);
	END GENERATE loop73;
	wire_rad_ff3c_w_q_range2365w(0) <= rad_ff3c(22);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff4c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff4c <= wire_alt_sqrt_block2_w_addnode_w4c_range237w;
			END IF;
		END IF;
	END PROCESS;
	loop74 : FOR i IN 0 TO 5 GENERATE 
		wire_rad_ff4c_w_lg_w_lg_w_q_range2397w2400w2401w(i) <= wire_rad_ff4c_w_lg_w_q_range2397w2400w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w5c_range2396w2399w(i);
	END GENERATE loop74;
	loop75 : FOR i IN 0 TO 5 GENERATE 
		wire_rad_ff4c_w_lg_w_q_range2397w2398w(i) <= wire_rad_ff4c_w_q_range2397w(0) AND wire_alt_sqrt_block2_w_qlevel_w5c_range2396w(i);
	END GENERATE loop75;
	wire_rad_ff4c_w_lg_w_q_range2397w2400w(0) <= NOT wire_rad_ff4c_w_q_range2397w(0);
	loop76 : FOR i IN 0 TO 5 GENERATE 
		wire_rad_ff4c_w_lg_w_lg_w_lg_w_q_range2397w2400w2401w2402w(i) <= wire_rad_ff4c_w_lg_w_lg_w_q_range2397w2400w2401w(i) OR wire_rad_ff4c_w_lg_w_q_range2397w2398w(i);
	END GENERATE loop76;
	wire_rad_ff4c_w_q_range2397w(0) <= rad_ff4c(21);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff5c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff5c <= wire_alt_sqrt_block2_w_addnode_w5c_range238w;
			END IF;
		END IF;
	END PROCESS;
	loop77 : FOR i IN 0 TO 6 GENERATE 
		wire_rad_ff5c_w_lg_w_lg_w_q_range2429w2432w2433w(i) <= wire_rad_ff5c_w_lg_w_q_range2429w2432w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w6c_range2428w2431w(i);
	END GENERATE loop77;
	loop78 : FOR i IN 0 TO 6 GENERATE 
		wire_rad_ff5c_w_lg_w_q_range2429w2430w(i) <= wire_rad_ff5c_w_q_range2429w(0) AND wire_alt_sqrt_block2_w_qlevel_w6c_range2428w(i);
	END GENERATE loop78;
	wire_rad_ff5c_w_lg_w_q_range2429w2432w(0) <= NOT wire_rad_ff5c_w_q_range2429w(0);
	loop79 : FOR i IN 0 TO 6 GENERATE 
		wire_rad_ff5c_w_lg_w_lg_w_lg_w_q_range2429w2432w2433w2434w(i) <= wire_rad_ff5c_w_lg_w_lg_w_q_range2429w2432w2433w(i) OR wire_rad_ff5c_w_lg_w_q_range2429w2430w(i);
	END GENERATE loop79;
	wire_rad_ff5c_w_q_range2429w(0) <= rad_ff5c(20);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff6c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff6c <= wire_alt_sqrt_block2_w_addnode_w6c_range239w;
			END IF;
		END IF;
	END PROCESS;
	loop80 : FOR i IN 0 TO 7 GENERATE 
		wire_rad_ff6c_w_lg_w_lg_w_q_range2461w2464w2465w(i) <= wire_rad_ff6c_w_lg_w_q_range2461w2464w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w7c_range2460w2463w(i);
	END GENERATE loop80;
	loop81 : FOR i IN 0 TO 7 GENERATE 
		wire_rad_ff6c_w_lg_w_q_range2461w2462w(i) <= wire_rad_ff6c_w_q_range2461w(0) AND wire_alt_sqrt_block2_w_qlevel_w7c_range2460w(i);
	END GENERATE loop81;
	wire_rad_ff6c_w_lg_w_q_range2461w2464w(0) <= NOT wire_rad_ff6c_w_q_range2461w(0);
	loop82 : FOR i IN 0 TO 7 GENERATE 
		wire_rad_ff6c_w_lg_w_lg_w_lg_w_q_range2461w2464w2465w2466w(i) <= wire_rad_ff6c_w_lg_w_lg_w_q_range2461w2464w2465w(i) OR wire_rad_ff6c_w_lg_w_q_range2461w2462w(i);
	END GENERATE loop82;
	wire_rad_ff6c_w_q_range2461w(0) <= rad_ff6c(19);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff7c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff7c <= wire_alt_sqrt_block2_w_addnode_w7c_range240w;
			END IF;
		END IF;
	END PROCESS;
	loop83 : FOR i IN 0 TO 8 GENERATE 
		wire_rad_ff7c_w_lg_w_lg_w_q_range2493w2496w2497w(i) <= wire_rad_ff7c_w_lg_w_q_range2493w2496w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w8c_range2492w2495w(i);
	END GENERATE loop83;
	loop84 : FOR i IN 0 TO 8 GENERATE 
		wire_rad_ff7c_w_lg_w_q_range2493w2494w(i) <= wire_rad_ff7c_w_q_range2493w(0) AND wire_alt_sqrt_block2_w_qlevel_w8c_range2492w(i);
	END GENERATE loop84;
	wire_rad_ff7c_w_lg_w_q_range2493w2496w(0) <= NOT wire_rad_ff7c_w_q_range2493w(0);
	loop85 : FOR i IN 0 TO 8 GENERATE 
		wire_rad_ff7c_w_lg_w_lg_w_lg_w_q_range2493w2496w2497w2498w(i) <= wire_rad_ff7c_w_lg_w_lg_w_q_range2493w2496w2497w(i) OR wire_rad_ff7c_w_lg_w_q_range2493w2494w(i);
	END GENERATE loop85;
	wire_rad_ff7c_w_q_range2493w(0) <= rad_ff7c(18);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff8c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff8c <= wire_alt_sqrt_block2_w_addnode_w8c_range241w;
			END IF;
		END IF;
	END PROCESS;
	loop86 : FOR i IN 0 TO 9 GENERATE 
		wire_rad_ff8c_w_lg_w_lg_w_q_range2525w2528w2529w(i) <= wire_rad_ff8c_w_lg_w_q_range2525w2528w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w9c_range2524w2527w(i);
	END GENERATE loop86;
	loop87 : FOR i IN 0 TO 9 GENERATE 
		wire_rad_ff8c_w_lg_w_q_range2525w2526w(i) <= wire_rad_ff8c_w_q_range2525w(0) AND wire_alt_sqrt_block2_w_qlevel_w9c_range2524w(i);
	END GENERATE loop87;
	wire_rad_ff8c_w_lg_w_q_range2525w2528w(0) <= NOT wire_rad_ff8c_w_q_range2525w(0);
	loop88 : FOR i IN 0 TO 9 GENERATE 
		wire_rad_ff8c_w_lg_w_lg_w_lg_w_q_range2525w2528w2529w2530w(i) <= wire_rad_ff8c_w_lg_w_lg_w_q_range2525w2528w2529w(i) OR wire_rad_ff8c_w_lg_w_q_range2525w2526w(i);
	END GENERATE loop88;
	wire_rad_ff8c_w_q_range2525w(0) <= rad_ff8c(17);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff9c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff9c <= wire_alt_sqrt_block2_w_addnode_w9c_range242w;
			END IF;
		END IF;
	END PROCESS;
	loop89 : FOR i IN 0 TO 10 GENERATE 
		wire_rad_ff9c_w_lg_w_lg_w_q_range2557w2560w2561w(i) <= wire_rad_ff9c_w_lg_w_q_range2557w2560w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w10c_range2556w2559w(i);
	END GENERATE loop89;
	loop90 : FOR i IN 0 TO 10 GENERATE 
		wire_rad_ff9c_w_lg_w_q_range2557w2558w(i) <= wire_rad_ff9c_w_q_range2557w(0) AND wire_alt_sqrt_block2_w_qlevel_w10c_range2556w(i);
	END GENERATE loop90;
	wire_rad_ff9c_w_lg_w_q_range2557w2560w(0) <= NOT wire_rad_ff9c_w_q_range2557w(0);
	loop91 : FOR i IN 0 TO 10 GENERATE 
		wire_rad_ff9c_w_lg_w_lg_w_lg_w_q_range2557w2560w2561w2562w(i) <= wire_rad_ff9c_w_lg_w_lg_w_q_range2557w2560w2561w(i) OR wire_rad_ff9c_w_lg_w_q_range2557w2558w(i);
	END GENERATE loop91;
	wire_rad_ff9c_w_q_range2557w(0) <= rad_ff9c(16);
	wire_add_sub10_dataa <= ( slevel_w6c(26 DOWNTO 18));
	wire_add_sub10_datab <= ( wire_rad_ff5c_w_lg_w_lg_w_lg_w_q_range2429w2432w2433w2434w & qlevel_w6c(1 DOWNTO 0));
	add_sub10 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => wire_add_sub10_dataa,
		datab => wire_add_sub10_datab,
		result => wire_add_sub10_result
	  );
	wire_add_sub11_dataa <= ( slevel_w7c(26 DOWNTO 17));
	wire_add_sub11_datab <= ( wire_rad_ff6c_w_lg_w_lg_w_lg_w_q_range2461w2464w2465w2466w & qlevel_w7c(1 DOWNTO 0));
	add_sub11 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 10
	  )
	  PORT MAP ( 
		dataa => wire_add_sub11_dataa,
		datab => wire_add_sub11_datab,
		result => wire_add_sub11_result
	  );
	wire_add_sub12_dataa <= ( slevel_w8c(26 DOWNTO 16));
	wire_add_sub12_datab <= ( wire_rad_ff7c_w_lg_w_lg_w_lg_w_q_range2493w2496w2497w2498w & qlevel_w8c(1 DOWNTO 0));
	add_sub12 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 11
	  )
	  PORT MAP ( 
		dataa => wire_add_sub12_dataa,
		datab => wire_add_sub12_datab,
		result => wire_add_sub12_result
	  );
	wire_add_sub13_dataa <= ( slevel_w9c(26 DOWNTO 15));
	wire_add_sub13_datab <= ( wire_rad_ff8c_w_lg_w_lg_w_lg_w_q_range2525w2528w2529w2530w & qlevel_w9c(1 DOWNTO 0));
	add_sub13 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 12
	  )
	  PORT MAP ( 
		dataa => wire_add_sub13_dataa,
		datab => wire_add_sub13_datab,
		result => wire_add_sub13_result
	  );
	wire_add_sub14_dataa <= ( slevel_w10c(26 DOWNTO 14));
	wire_add_sub14_datab <= ( wire_rad_ff9c_w_lg_w_lg_w_lg_w_q_range2557w2560w2561w2562w & qlevel_w10c(1 DOWNTO 0));
	add_sub14 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		dataa => wire_add_sub14_dataa,
		datab => wire_add_sub14_datab,
		result => wire_add_sub14_result
	  );
	wire_add_sub15_dataa <= ( slevel_w11c(26 DOWNTO 13));
	wire_add_sub15_datab <= ( wire_rad_ff10c_w_lg_w_lg_w_lg_w_q_range2589w2592w2593w2594w & qlevel_w11c(1 DOWNTO 0));
	add_sub15 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 14
	  )
	  PORT MAP ( 
		dataa => wire_add_sub15_dataa,
		datab => wire_add_sub15_datab,
		result => wire_add_sub15_result
	  );
	wire_add_sub16_dataa <= ( slevel_w12c(26 DOWNTO 13));
	wire_add_sub16_datab <= ( wire_rad_ff11c_w_lg_w_lg_w_lg_w_q_range2620w2623w2624w2625w & qlevel_w12c(1));
	add_sub16 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 14
	  )
	  PORT MAP ( 
		dataa => wire_add_sub16_dataa,
		datab => wire_add_sub16_datab,
		result => wire_add_sub16_result
	  );
	wire_add_sub17_dataa <= ( slevel_w13c(26 DOWNTO 14));
	wire_add_sub17_datab <= ( wire_rad_ff12c_w_lg_w_lg_w_lg_w_q_range2652w2655w2656w2657w);
	add_sub17 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		dataa => wire_add_sub17_dataa,
		datab => wire_add_sub17_datab,
		result => wire_add_sub17_result
	  );
	wire_add_sub18_dataa <= ( slevel_w14c(26 DOWNTO 13));
	wire_add_sub18_datab <= ( wire_rad_ff13c_w_lg_w_lg_w_lg_w_q_range2691w2694w2695w2696w);
	add_sub18 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 14
	  )
	  PORT MAP ( 
		dataa => wire_add_sub18_dataa,
		datab => wire_add_sub18_datab,
		result => wire_add_sub18_result
	  );
	wire_add_sub19_dataa <= ( slevel_w15c(26 DOWNTO 12));
	wire_add_sub19_datab <= ( wire_rad_ff14c_w_lg_w_lg_w_lg_w_q_range2730w2733w2734w2735w);
	add_sub19 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 15
	  )
	  PORT MAP ( 
		dataa => wire_add_sub19_dataa,
		datab => wire_add_sub19_datab,
		result => wire_add_sub19_result
	  );
	wire_add_sub20_dataa <= ( slevel_w16c(26 DOWNTO 11));
	wire_add_sub20_datab <= ( wire_rad_ff15c_w_lg_w_lg_w_lg_w_q_range2769w2772w2773w2774w);
	add_sub20 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 16
	  )
	  PORT MAP ( 
		dataa => wire_add_sub20_dataa,
		datab => wire_add_sub20_datab,
		result => wire_add_sub20_result
	  );
	wire_add_sub21_dataa <= ( slevel_w17c(26 DOWNTO 10));
	wire_add_sub21_datab <= ( wire_rad_ff16c_w_lg_w_lg_w_lg_w_q_range2808w2811w2812w2813w);
	add_sub21 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 17
	  )
	  PORT MAP ( 
		dataa => wire_add_sub21_dataa,
		datab => wire_add_sub21_datab,
		result => wire_add_sub21_result
	  );
	wire_add_sub22_dataa <= ( slevel_w18c(26 DOWNTO 9));
	wire_add_sub22_datab <= ( wire_rad_ff17c_w_lg_w_lg_w_lg_w_q_range2847w2850w2851w2852w);
	add_sub22 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 18
	  )
	  PORT MAP ( 
		dataa => wire_add_sub22_dataa,
		datab => wire_add_sub22_datab,
		result => wire_add_sub22_result
	  );
	wire_add_sub23_dataa <= ( slevel_w19c(26 DOWNTO 8));
	wire_add_sub23_datab <= ( wire_rad_ff18c_w_lg_w_lg_w_lg_w_q_range2886w2889w2890w2891w);
	add_sub23 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 19
	  )
	  PORT MAP ( 
		dataa => wire_add_sub23_dataa,
		datab => wire_add_sub23_datab,
		result => wire_add_sub23_result
	  );
	wire_add_sub24_dataa <= ( slevel_w20c(26 DOWNTO 7));
	wire_add_sub24_datab <= ( wire_rad_ff19c_w_lg_w_lg_w_lg_w_q_range2925w2928w2929w2930w);
	add_sub24 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 20
	  )
	  PORT MAP ( 
		dataa => wire_add_sub24_dataa,
		datab => wire_add_sub24_datab,
		result => wire_add_sub24_result
	  );
	wire_add_sub25_dataa <= ( slevel_w21c(26 DOWNTO 6));
	wire_add_sub25_datab <= ( wire_rad_ff20c_w_lg_w_lg_w_lg_w_q_range2964w2967w2968w2969w);
	add_sub25 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 21
	  )
	  PORT MAP ( 
		dataa => wire_add_sub25_dataa,
		datab => wire_add_sub25_datab,
		result => wire_add_sub25_result
	  );
	wire_add_sub26_dataa <= ( slevel_w22c(26 DOWNTO 5));
	wire_add_sub26_datab <= ( wire_rad_ff21c_w_lg_w_lg_w_lg_w_q_range3003w3006w3007w3008w);
	add_sub26 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 22
	  )
	  PORT MAP ( 
		dataa => wire_add_sub26_dataa,
		datab => wire_add_sub26_datab,
		result => wire_add_sub26_result
	  );
	wire_add_sub27_dataa <= ( slevel_w23c(26 DOWNTO 4));
	wire_add_sub27_datab <= ( wire_rad_ff22c_w_lg_w_lg_w_lg_w_q_range3042w3045w3046w3047w);
	add_sub27 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 23
	  )
	  PORT MAP ( 
		dataa => wire_add_sub27_dataa,
		datab => wire_add_sub27_datab,
		result => wire_add_sub27_result
	  );
	wire_add_sub28_dataa <= ( slevel_w24c(26 DOWNTO 3));
	wire_add_sub28_datab <= ( qlevel_w24c(26 DOWNTO 25) & wire_rad_ff23c_w_lg_w_lg_w_lg_w_q_range3069w3070w3086w3087w);
	add_sub28 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 24
	  )
	  PORT MAP ( 
		dataa => wire_add_sub28_dataa,
		datab => wire_add_sub28_datab,
		result => wire_add_sub28_result
	  );
	wire_add_sub4_dataa <= ( slevel_w0c(26 DOWNTO 24));
	wire_add_sub4_datab <= ( qlevel_w0c(2 DOWNTO 0));
	add_sub4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 3
	  )
	  PORT MAP ( 
		dataa => wire_add_sub4_dataa,
		datab => wire_add_sub4_datab,
		result => wire_add_sub4_result
	  );
	wire_add_sub5_dataa <= ( slevel_w1c(26 DOWNTO 23));
	wire_add_sub5_datab <= ( qlevel_w1c(3 DOWNTO 0));
	add_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		dataa => wire_add_sub5_dataa,
		datab => wire_add_sub5_datab,
		result => wire_add_sub5_result
	  );
	wire_add_sub6_dataa <= ( slevel_w2c(26 DOWNTO 22));
	wire_add_sub6_datab <= ( wire_rad_ff1c_w_lg_w_lg_w_lg_w_q_range2301w2304w2305w2306w & qlevel_w2c(1 DOWNTO 0));
	add_sub6 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		dataa => wire_add_sub6_dataa,
		datab => wire_add_sub6_datab,
		result => wire_add_sub6_result
	  );
	wire_add_sub7_dataa <= ( slevel_w3c(26 DOWNTO 21));
	wire_add_sub7_datab <= ( wire_rad_ff2c_w_lg_w_lg_w_lg_w_q_range2333w2336w2337w2338w & qlevel_w3c(1 DOWNTO 0));
	add_sub7 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		dataa => wire_add_sub7_dataa,
		datab => wire_add_sub7_datab,
		result => wire_add_sub7_result
	  );
	wire_add_sub8_dataa <= ( slevel_w4c(26 DOWNTO 20));
	wire_add_sub8_datab <= ( wire_rad_ff3c_w_lg_w_lg_w_lg_w_q_range2365w2368w2369w2370w & qlevel_w4c(1 DOWNTO 0));
	add_sub8 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 7
	  )
	  PORT MAP ( 
		dataa => wire_add_sub8_dataa,
		datab => wire_add_sub8_datab,
		result => wire_add_sub8_result
	  );
	wire_add_sub9_dataa <= ( slevel_w5c(26 DOWNTO 19));
	wire_add_sub9_datab <= ( wire_rad_ff4c_w_lg_w_lg_w_lg_w_q_range2397w2400w2401w2402w & qlevel_w5c(1 DOWNTO 0));
	add_sub9 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		dataa => wire_add_sub9_dataa,
		datab => wire_add_sub9_datab,
		result => wire_add_sub9_result
	  );

 END RTL; --k_ukf_sqrt_alt_sqrt_block_nfb

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 27 reg 1433 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  k_ukf_sqrt_altfp_sqrt_0mc IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END k_ukf_sqrt_altfp_sqrt_0mc;

 ARCHITECTURE RTL OF k_ukf_sqrt_altfp_sqrt_0mc IS

	 SIGNAL  wire_alt_sqrt_block2_root_result	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL	 exp_all_one_ff	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff1	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff20c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff210c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff211c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff212c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff213c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff214c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff215c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff216c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff217c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff218c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff219c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff21c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff220c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff221c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff222c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff223c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff224c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff22c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff23c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff24c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff25c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff26c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff27c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff28c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff29c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_in_ff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range27w31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range32w36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range37w41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range42w46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range47w51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range52w56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range57w61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range27w29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range32w34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range37w39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range42w44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range47w49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range52w54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range57w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exp_not_zero_ff	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_ff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff23	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff24	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_in_ff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range62w159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range161w162w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range163w164w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range128w168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_lg_w_q_range163w164w165w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range92w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range95w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range98w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range101w103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range104w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range107w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range110w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range113w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range116w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range119w121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range65w67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range122w124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range125w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range128w130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range68w70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range71w73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range74w76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range77w79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range80w82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range83w85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range86w88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range89w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range161w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range163w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 man_not_zero_ff	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_not_zero_ff_w_lg_q131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 man_result_ff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_rounding_ff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_rounding_ff_w_lg_q177w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_man_rounding_ff_w_lg_w_lg_q177w178w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL	 nan_man_ff0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff23	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff24	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_sign_node_ff_w_lg_q136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 sign_node_ff2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff23	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff24	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff25	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff26	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff27	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff23	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff24	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_sub1_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub1_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub3_datab	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_add_sub3_result	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_ff2_w152w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_preadjust_w160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exp_ff2_w152w153w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_exp_ff2_w152w153w154w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_preadjust_w169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  bias :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  exp_all_one_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_div_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_ff2_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_not_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  infinitycondition_w :	STD_LOGIC;
	 SIGNAL  man_not_zero_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_root_result_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  nancondition_w :	STD_LOGIC;
	 SIGNAL  preadjust_w :	STD_LOGIC;
	 SIGNAL  radicand_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  roundbit_w :	STD_LOGIC;
	 SIGNAL  wire_w_data_range21w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_data_range20w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  k_ukf_sqrt_alt_sqrt_block_nfb
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		rad	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0);
		root_result	:	OUT  STD_LOGIC_VECTOR(24 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	loop92 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_exp_ff2_w152w(i) <= exp_ff2_w(i) AND zero_exp_ff24;
	END GENERATE loop92;
	wire_w_lg_preadjust_w160w(0) <= NOT preadjust_w;
	loop93 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_exp_ff2_w152w153w(i) <= wire_w_lg_exp_ff2_w152w(i) OR nan_man_ff24;
	END GENERATE loop93;
	loop94 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_w_lg_exp_ff2_w152w153w154w(i) <= wire_w_lg_w_lg_exp_ff2_w152w153w(i) OR infinity_ff24;
	END GENERATE loop94;
	wire_w_lg_preadjust_w169w(0) <= preadjust_w OR wire_man_in_ff_w_lg_w_q_range128w168w(0);
	aclr <= '0';
	bias <= ( "0" & "1" & "1" & "1" & "1" & "1" & "1" & "1");
	clk_en <= '1';
	exp_all_one_w <= ( wire_exp_in_ff_w_lg_w_q_range57w61w & wire_exp_in_ff_w_lg_w_q_range52w56w & wire_exp_in_ff_w_lg_w_q_range47w51w & wire_exp_in_ff_w_lg_w_q_range42w46w & wire_exp_in_ff_w_lg_w_q_range37w41w & wire_exp_in_ff_w_lg_w_q_range32w36w & wire_exp_in_ff_w_lg_w_q_range27w31w & exp_in_ff(0));
	exp_div_w <= ( wire_add_sub1_result(8 DOWNTO 1));
	exp_ff2_w <= exp_ff224c;
	exp_not_zero_w <= ( wire_exp_in_ff_w_lg_w_q_range57w59w & wire_exp_in_ff_w_lg_w_q_range52w54w & wire_exp_in_ff_w_lg_w_q_range47w49w & wire_exp_in_ff_w_lg_w_q_range42w44w & wire_exp_in_ff_w_lg_w_q_range37w39w & wire_exp_in_ff_w_lg_w_q_range32w34w & wire_exp_in_ff_w_lg_w_q_range27w29w & exp_in_ff(0));
	infinitycondition_w <= (wire_man_not_zero_ff_w_lg_q131w(0) AND exp_all_one_ff);
	man_not_zero_w <= ( wire_man_in_ff_w_lg_w_q_range128w130w & wire_man_in_ff_w_lg_w_q_range125w127w & wire_man_in_ff_w_lg_w_q_range122w124w & wire_man_in_ff_w_lg_w_q_range119w121w & wire_man_in_ff_w_lg_w_q_range116w118w & wire_man_in_ff_w_lg_w_q_range113w115w & wire_man_in_ff_w_lg_w_q_range110w112w & wire_man_in_ff_w_lg_w_q_range107w109w & wire_man_in_ff_w_lg_w_q_range104w106w & wire_man_in_ff_w_lg_w_q_range101w103w & wire_man_in_ff_w_lg_w_q_range98w100w & wire_man_in_ff_w_lg_w_q_range95w97w & wire_man_in_ff_w_lg_w_q_range92w94w & wire_man_in_ff_w_lg_w_q_range89w91w & wire_man_in_ff_w_lg_w_q_range86w88w & wire_man_in_ff_w_lg_w_q_range83w85w & wire_man_in_ff_w_lg_w_q_range80w82w & wire_man_in_ff_w_lg_w_q_range77w79w & wire_man_in_ff_w_lg_w_q_range74w76w & wire_man_in_ff_w_lg_w_q_range71w73w & wire_man_in_ff_w_lg_w_q_range68w70w & wire_man_in_ff_w_lg_w_q_range65w67w & man_in_ff(0));
	man_root_result_w <= wire_alt_sqrt_block2_root_result;
	nancondition_w <= ((sign_node_ff1 AND exp_not_zero_ff) OR (exp_all_one_ff AND man_not_zero_ff));
	preadjust_w <= exp_in_ff(0);
	radicand_w <= ( wire_w_lg_preadjust_w160w & wire_w_lg_preadjust_w169w & wire_man_in_ff_w_lg_w_lg_w_q_range163w164w165w & wire_man_in_ff_w_lg_w_q_range62w159w & "0");
	result <= ( sign_node_ff27 & exp_result_ff & man_result_ff);
	roundbit_w <= wire_alt_sqrt_block2_root_result(0);
	wire_w_data_range21w <= data(22 DOWNTO 0);
	wire_w_data_range20w <= data(30 DOWNTO 23);
	wire_w_exp_all_one_w_range25w(0) <= exp_all_one_w(0);
	wire_w_exp_all_one_w_range30w(0) <= exp_all_one_w(1);
	wire_w_exp_all_one_w_range35w(0) <= exp_all_one_w(2);
	wire_w_exp_all_one_w_range40w(0) <= exp_all_one_w(3);
	wire_w_exp_all_one_w_range45w(0) <= exp_all_one_w(4);
	wire_w_exp_all_one_w_range50w(0) <= exp_all_one_w(5);
	wire_w_exp_all_one_w_range55w(0) <= exp_all_one_w(6);
	wire_w_exp_not_zero_w_range23w(0) <= exp_not_zero_w(0);
	wire_w_exp_not_zero_w_range28w(0) <= exp_not_zero_w(1);
	wire_w_exp_not_zero_w_range33w(0) <= exp_not_zero_w(2);
	wire_w_exp_not_zero_w_range38w(0) <= exp_not_zero_w(3);
	wire_w_exp_not_zero_w_range43w(0) <= exp_not_zero_w(4);
	wire_w_exp_not_zero_w_range48w(0) <= exp_not_zero_w(5);
	wire_w_exp_not_zero_w_range53w(0) <= exp_not_zero_w(6);
	wire_w_man_not_zero_w_range63w(0) <= man_not_zero_w(0);
	wire_w_man_not_zero_w_range93w(0) <= man_not_zero_w(10);
	wire_w_man_not_zero_w_range96w(0) <= man_not_zero_w(11);
	wire_w_man_not_zero_w_range99w(0) <= man_not_zero_w(12);
	wire_w_man_not_zero_w_range102w(0) <= man_not_zero_w(13);
	wire_w_man_not_zero_w_range105w(0) <= man_not_zero_w(14);
	wire_w_man_not_zero_w_range108w(0) <= man_not_zero_w(15);
	wire_w_man_not_zero_w_range111w(0) <= man_not_zero_w(16);
	wire_w_man_not_zero_w_range114w(0) <= man_not_zero_w(17);
	wire_w_man_not_zero_w_range117w(0) <= man_not_zero_w(18);
	wire_w_man_not_zero_w_range120w(0) <= man_not_zero_w(19);
	wire_w_man_not_zero_w_range66w(0) <= man_not_zero_w(1);
	wire_w_man_not_zero_w_range123w(0) <= man_not_zero_w(20);
	wire_w_man_not_zero_w_range126w(0) <= man_not_zero_w(21);
	wire_w_man_not_zero_w_range69w(0) <= man_not_zero_w(2);
	wire_w_man_not_zero_w_range72w(0) <= man_not_zero_w(3);
	wire_w_man_not_zero_w_range75w(0) <= man_not_zero_w(4);
	wire_w_man_not_zero_w_range78w(0) <= man_not_zero_w(5);
	wire_w_man_not_zero_w_range81w(0) <= man_not_zero_w(6);
	wire_w_man_not_zero_w_range84w(0) <= man_not_zero_w(7);
	wire_w_man_not_zero_w_range87w(0) <= man_not_zero_w(8);
	wire_w_man_not_zero_w_range90w(0) <= man_not_zero_w(9);
	alt_sqrt_block2 :  k_ukf_sqrt_alt_sqrt_block_nfb
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		rad => radicand_w,
		root_result => wire_alt_sqrt_block2_root_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_all_one_ff <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_all_one_ff <= exp_all_one_w(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff1 <= exp_div_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff20c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff20c <= exp_ff1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff210c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff210c <= exp_ff29c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff211c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff211c <= exp_ff210c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff212c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff212c <= exp_ff211c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff213c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff213c <= exp_ff212c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff214c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff214c <= exp_ff213c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff215c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff215c <= exp_ff214c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff216c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff216c <= exp_ff215c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff217c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff217c <= exp_ff216c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff218c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff218c <= exp_ff217c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff219c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff219c <= exp_ff218c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff21c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff21c <= exp_ff20c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff220c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff220c <= exp_ff219c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff221c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff221c <= exp_ff220c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff222c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff222c <= exp_ff221c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff223c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff223c <= exp_ff222c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff224c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff224c <= exp_ff223c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff22c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff22c <= exp_ff21c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff23c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff23c <= exp_ff22c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff24c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff24c <= exp_ff23c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff25c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff25c <= exp_ff24c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff26c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff26c <= exp_ff25c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff27c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff27c <= exp_ff26c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff28c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff28c <= exp_ff27c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff29c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff29c <= exp_ff28c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_in_ff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_in_ff <= wire_w_data_range20w;
			END IF;
		END IF;
	END PROCESS;
	wire_exp_in_ff_w_lg_w_q_range27w31w(0) <= wire_exp_in_ff_w_q_range27w(0) AND wire_w_exp_all_one_w_range25w(0);
	wire_exp_in_ff_w_lg_w_q_range32w36w(0) <= wire_exp_in_ff_w_q_range32w(0) AND wire_w_exp_all_one_w_range30w(0);
	wire_exp_in_ff_w_lg_w_q_range37w41w(0) <= wire_exp_in_ff_w_q_range37w(0) AND wire_w_exp_all_one_w_range35w(0);
	wire_exp_in_ff_w_lg_w_q_range42w46w(0) <= wire_exp_in_ff_w_q_range42w(0) AND wire_w_exp_all_one_w_range40w(0);
	wire_exp_in_ff_w_lg_w_q_range47w51w(0) <= wire_exp_in_ff_w_q_range47w(0) AND wire_w_exp_all_one_w_range45w(0);
	wire_exp_in_ff_w_lg_w_q_range52w56w(0) <= wire_exp_in_ff_w_q_range52w(0) AND wire_w_exp_all_one_w_range50w(0);
	wire_exp_in_ff_w_lg_w_q_range57w61w(0) <= wire_exp_in_ff_w_q_range57w(0) AND wire_w_exp_all_one_w_range55w(0);
	wire_exp_in_ff_w_lg_w_q_range27w29w(0) <= wire_exp_in_ff_w_q_range27w(0) OR wire_w_exp_not_zero_w_range23w(0);
	wire_exp_in_ff_w_lg_w_q_range32w34w(0) <= wire_exp_in_ff_w_q_range32w(0) OR wire_w_exp_not_zero_w_range28w(0);
	wire_exp_in_ff_w_lg_w_q_range37w39w(0) <= wire_exp_in_ff_w_q_range37w(0) OR wire_w_exp_not_zero_w_range33w(0);
	wire_exp_in_ff_w_lg_w_q_range42w44w(0) <= wire_exp_in_ff_w_q_range42w(0) OR wire_w_exp_not_zero_w_range38w(0);
	wire_exp_in_ff_w_lg_w_q_range47w49w(0) <= wire_exp_in_ff_w_q_range47w(0) OR wire_w_exp_not_zero_w_range43w(0);
	wire_exp_in_ff_w_lg_w_q_range52w54w(0) <= wire_exp_in_ff_w_q_range52w(0) OR wire_w_exp_not_zero_w_range48w(0);
	wire_exp_in_ff_w_lg_w_q_range57w59w(0) <= wire_exp_in_ff_w_q_range57w(0) OR wire_w_exp_not_zero_w_range53w(0);
	wire_exp_in_ff_w_q_range27w(0) <= exp_in_ff(1);
	wire_exp_in_ff_w_q_range32w(0) <= exp_in_ff(2);
	wire_exp_in_ff_w_q_range37w(0) <= exp_in_ff(3);
	wire_exp_in_ff_w_q_range42w(0) <= exp_in_ff(4);
	wire_exp_in_ff_w_q_range47w(0) <= exp_in_ff(5);
	wire_exp_in_ff_w_q_range52w(0) <= exp_in_ff(6);
	wire_exp_in_ff_w_q_range57w(0) <= exp_in_ff(7);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_not_zero_ff <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_not_zero_ff <= exp_not_zero_w(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_ff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_ff <= wire_w_lg_w_lg_w_lg_exp_ff2_w152w153w154w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff0 <= (infinitycondition_w AND wire_sign_node_ff_w_lg_q136w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff1 <= infinity_ff0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff2 <= infinity_ff1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff3 <= infinity_ff2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff4 <= infinity_ff3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff5 <= infinity_ff4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff6 <= infinity_ff5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff7 <= infinity_ff6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff8 <= infinity_ff7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff9 <= infinity_ff8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff10 <= infinity_ff9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff11 <= infinity_ff10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff12 <= infinity_ff11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff13 <= infinity_ff12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff14 <= infinity_ff13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff15 <= infinity_ff14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff16 <= infinity_ff15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff17 <= infinity_ff16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff18 <= infinity_ff17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff19 <= infinity_ff18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff20 <= infinity_ff19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff21 <= infinity_ff20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff22 <= infinity_ff21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff23 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff23 <= infinity_ff22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff24 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff24 <= infinity_ff23;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_in_ff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_in_ff <= wire_w_data_range21w;
			END IF;
		END IF;
	END PROCESS;
	wire_man_in_ff_w_lg_w_q_range62w159w(0) <= wire_man_in_ff_w_q_range62w(0) AND preadjust_w;
	loop95 : FOR i IN 0 TO 21 GENERATE 
		wire_man_in_ff_w_lg_w_q_range161w162w(i) <= wire_man_in_ff_w_q_range161w(i) AND wire_w_lg_preadjust_w160w(0);
	END GENERATE loop95;
	loop96 : FOR i IN 0 TO 21 GENERATE 
		wire_man_in_ff_w_lg_w_q_range163w164w(i) <= wire_man_in_ff_w_q_range163w(i) AND preadjust_w;
	END GENERATE loop96;
	wire_man_in_ff_w_lg_w_q_range128w168w(0) <= wire_man_in_ff_w_q_range128w(0) AND wire_w_lg_preadjust_w160w(0);
	loop97 : FOR i IN 0 TO 21 GENERATE 
		wire_man_in_ff_w_lg_w_lg_w_q_range163w164w165w(i) <= wire_man_in_ff_w_lg_w_q_range163w164w(i) OR wire_man_in_ff_w_lg_w_q_range161w162w(i);
	END GENERATE loop97;
	wire_man_in_ff_w_lg_w_q_range92w94w(0) <= wire_man_in_ff_w_q_range92w(0) OR wire_w_man_not_zero_w_range90w(0);
	wire_man_in_ff_w_lg_w_q_range95w97w(0) <= wire_man_in_ff_w_q_range95w(0) OR wire_w_man_not_zero_w_range93w(0);
	wire_man_in_ff_w_lg_w_q_range98w100w(0) <= wire_man_in_ff_w_q_range98w(0) OR wire_w_man_not_zero_w_range96w(0);
	wire_man_in_ff_w_lg_w_q_range101w103w(0) <= wire_man_in_ff_w_q_range101w(0) OR wire_w_man_not_zero_w_range99w(0);
	wire_man_in_ff_w_lg_w_q_range104w106w(0) <= wire_man_in_ff_w_q_range104w(0) OR wire_w_man_not_zero_w_range102w(0);
	wire_man_in_ff_w_lg_w_q_range107w109w(0) <= wire_man_in_ff_w_q_range107w(0) OR wire_w_man_not_zero_w_range105w(0);
	wire_man_in_ff_w_lg_w_q_range110w112w(0) <= wire_man_in_ff_w_q_range110w(0) OR wire_w_man_not_zero_w_range108w(0);
	wire_man_in_ff_w_lg_w_q_range113w115w(0) <= wire_man_in_ff_w_q_range113w(0) OR wire_w_man_not_zero_w_range111w(0);
	wire_man_in_ff_w_lg_w_q_range116w118w(0) <= wire_man_in_ff_w_q_range116w(0) OR wire_w_man_not_zero_w_range114w(0);
	wire_man_in_ff_w_lg_w_q_range119w121w(0) <= wire_man_in_ff_w_q_range119w(0) OR wire_w_man_not_zero_w_range117w(0);
	wire_man_in_ff_w_lg_w_q_range65w67w(0) <= wire_man_in_ff_w_q_range65w(0) OR wire_w_man_not_zero_w_range63w(0);
	wire_man_in_ff_w_lg_w_q_range122w124w(0) <= wire_man_in_ff_w_q_range122w(0) OR wire_w_man_not_zero_w_range120w(0);
	wire_man_in_ff_w_lg_w_q_range125w127w(0) <= wire_man_in_ff_w_q_range125w(0) OR wire_w_man_not_zero_w_range123w(0);
	wire_man_in_ff_w_lg_w_q_range128w130w(0) <= wire_man_in_ff_w_q_range128w(0) OR wire_w_man_not_zero_w_range126w(0);
	wire_man_in_ff_w_lg_w_q_range68w70w(0) <= wire_man_in_ff_w_q_range68w(0) OR wire_w_man_not_zero_w_range66w(0);
	wire_man_in_ff_w_lg_w_q_range71w73w(0) <= wire_man_in_ff_w_q_range71w(0) OR wire_w_man_not_zero_w_range69w(0);
	wire_man_in_ff_w_lg_w_q_range74w76w(0) <= wire_man_in_ff_w_q_range74w(0) OR wire_w_man_not_zero_w_range72w(0);
	wire_man_in_ff_w_lg_w_q_range77w79w(0) <= wire_man_in_ff_w_q_range77w(0) OR wire_w_man_not_zero_w_range75w(0);
	wire_man_in_ff_w_lg_w_q_range80w82w(0) <= wire_man_in_ff_w_q_range80w(0) OR wire_w_man_not_zero_w_range78w(0);
	wire_man_in_ff_w_lg_w_q_range83w85w(0) <= wire_man_in_ff_w_q_range83w(0) OR wire_w_man_not_zero_w_range81w(0);
	wire_man_in_ff_w_lg_w_q_range86w88w(0) <= wire_man_in_ff_w_q_range86w(0) OR wire_w_man_not_zero_w_range84w(0);
	wire_man_in_ff_w_lg_w_q_range89w91w(0) <= wire_man_in_ff_w_q_range89w(0) OR wire_w_man_not_zero_w_range87w(0);
	wire_man_in_ff_w_q_range62w(0) <= man_in_ff(0);
	wire_man_in_ff_w_q_range92w(0) <= man_in_ff(10);
	wire_man_in_ff_w_q_range95w(0) <= man_in_ff(11);
	wire_man_in_ff_w_q_range98w(0) <= man_in_ff(12);
	wire_man_in_ff_w_q_range101w(0) <= man_in_ff(13);
	wire_man_in_ff_w_q_range104w(0) <= man_in_ff(14);
	wire_man_in_ff_w_q_range107w(0) <= man_in_ff(15);
	wire_man_in_ff_w_q_range110w(0) <= man_in_ff(16);
	wire_man_in_ff_w_q_range113w(0) <= man_in_ff(17);
	wire_man_in_ff_w_q_range116w(0) <= man_in_ff(18);
	wire_man_in_ff_w_q_range119w(0) <= man_in_ff(19);
	wire_man_in_ff_w_q_range65w(0) <= man_in_ff(1);
	wire_man_in_ff_w_q_range122w(0) <= man_in_ff(20);
	wire_man_in_ff_w_q_range161w <= man_in_ff(21 DOWNTO 0);
	wire_man_in_ff_w_q_range125w(0) <= man_in_ff(21);
	wire_man_in_ff_w_q_range163w <= man_in_ff(22 DOWNTO 1);
	wire_man_in_ff_w_q_range128w(0) <= man_in_ff(22);
	wire_man_in_ff_w_q_range68w(0) <= man_in_ff(2);
	wire_man_in_ff_w_q_range71w(0) <= man_in_ff(3);
	wire_man_in_ff_w_q_range74w(0) <= man_in_ff(4);
	wire_man_in_ff_w_q_range77w(0) <= man_in_ff(5);
	wire_man_in_ff_w_q_range80w(0) <= man_in_ff(6);
	wire_man_in_ff_w_q_range83w(0) <= man_in_ff(7);
	wire_man_in_ff_w_q_range86w(0) <= man_in_ff(8);
	wire_man_in_ff_w_q_range89w(0) <= man_in_ff(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_not_zero_ff <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_not_zero_ff <= man_not_zero_w(22);
			END IF;
		END IF;
	END PROCESS;
	wire_man_not_zero_ff_w_lg_q131w(0) <= NOT man_not_zero_ff;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_result_ff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_result_ff <= wire_man_rounding_ff_w_lg_w_lg_q177w178w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_rounding_ff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_rounding_ff <= wire_add_sub3_result;
			END IF;
		END IF;
	END PROCESS;
	loop98 : FOR i IN 0 TO 22 GENERATE 
		wire_man_rounding_ff_w_lg_q177w(i) <= man_rounding_ff(i) AND zero_exp_ff24;
	END GENERATE loop98;
	loop99 : FOR i IN 0 TO 22 GENERATE 
		wire_man_rounding_ff_w_lg_w_lg_q177w178w(i) <= wire_man_rounding_ff_w_lg_q177w(i) OR nan_man_ff24;
	END GENERATE loop99;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff0 <= nancondition_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff1 <= nan_man_ff0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff2 <= nan_man_ff1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff3 <= nan_man_ff2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff4 <= nan_man_ff3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff5 <= nan_man_ff4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff6 <= nan_man_ff5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff7 <= nan_man_ff6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff8 <= nan_man_ff7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff9 <= nan_man_ff8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff10 <= nan_man_ff9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff11 <= nan_man_ff10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff12 <= nan_man_ff11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff13 <= nan_man_ff12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff14 <= nan_man_ff13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff15 <= nan_man_ff14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff16 <= nan_man_ff15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff17 <= nan_man_ff16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff18 <= nan_man_ff17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff19 <= nan_man_ff18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff20 <= nan_man_ff19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff21 <= nan_man_ff20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff22 <= nan_man_ff21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff23 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff23 <= nan_man_ff22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff24 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff24 <= nan_man_ff23;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff0 <= data(31);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff1 <= sign_node_ff0;
			END IF;
		END IF;
	END PROCESS;
	wire_sign_node_ff_w_lg_q136w(0) <= NOT sign_node_ff1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff2 <= sign_node_ff1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff3 <= sign_node_ff2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff4 <= sign_node_ff3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff5 <= sign_node_ff4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff6 <= sign_node_ff5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff7 <= sign_node_ff6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff8 <= sign_node_ff7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff9 <= sign_node_ff8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff10 <= sign_node_ff9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff11 <= sign_node_ff10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff12 <= sign_node_ff11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff13 <= sign_node_ff12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff14 <= sign_node_ff13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff15 <= sign_node_ff14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff16 <= sign_node_ff15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff17 <= sign_node_ff16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff18 <= sign_node_ff17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff19 <= sign_node_ff18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff20 <= sign_node_ff19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff21 <= sign_node_ff20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff22 <= sign_node_ff21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff23 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff23 <= sign_node_ff22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff24 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff24 <= sign_node_ff23;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff25 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff25 <= sign_node_ff24;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff26 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff26 <= sign_node_ff25;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff27 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff27 <= sign_node_ff26;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff0 <= exp_not_zero_ff;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff1 <= zero_exp_ff0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff2 <= zero_exp_ff1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff3 <= zero_exp_ff2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff4 <= zero_exp_ff3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff5 <= zero_exp_ff4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff6 <= zero_exp_ff5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff7 <= zero_exp_ff6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff8 <= zero_exp_ff7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff9 <= zero_exp_ff8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff10 <= zero_exp_ff9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff11 <= zero_exp_ff10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff12 <= zero_exp_ff11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff13 <= zero_exp_ff12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff14 <= zero_exp_ff13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff15 <= zero_exp_ff14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff16 <= zero_exp_ff15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff17 <= zero_exp_ff16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff18 <= zero_exp_ff17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff19 <= zero_exp_ff18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff20 <= zero_exp_ff19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff21 <= zero_exp_ff20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff22 <= zero_exp_ff21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff23 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff23 <= zero_exp_ff22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff24 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff24 <= zero_exp_ff23;
			END IF;
		END IF;
	END PROCESS;
	wire_add_sub1_dataa <= ( "0" & exp_in_ff);
	wire_add_sub1_datab <= ( "0" & bias);
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => wire_add_sub1_dataa,
		datab => wire_add_sub1_datab,
		result => wire_add_sub1_result
	  );
	wire_add_sub3_datab <= ( "0000000000000000000000" & roundbit_w);
	add_sub3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 23
	  )
	  PORT MAP ( 
		dataa => man_root_result_w(23 DOWNTO 1),
		datab => wire_add_sub3_datab,
		result => wire_add_sub3_result
	  );

 END RTL; --k_ukf_sqrt_altfp_sqrt_0mc
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY k_ukf_sqrt IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END k_ukf_sqrt;


ARCHITECTURE RTL OF k_ukf_sqrt IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT k_ukf_sqrt_altfp_sqrt_0mc
	PORT (
			clock	: IN STD_LOGIC ;
			data	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	k_ukf_sqrt_altfp_sqrt_0mc_component : k_ukf_sqrt_altfp_sqrt_0mc
	PORT MAP (
		clock => clock,
		data => data,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: FPM_FORMAT NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "1"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "28"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: data 0 0 32 0 INPUT NODEFVAL "data[31..0]"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data 0 0 32 0 data 0 0 32 0
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL k_ukf_sqrt.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL k_ukf_sqrt.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL k_ukf_sqrt.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL k_ukf_sqrt.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL k_ukf_sqrt_inst.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL k_ukf_sqrt_syn.v TRUE
-- Retrieval info: LIB_FILE: lpm
